library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.Types.all;

package Layer1_Weights is
constant weight_matrix_layer1 :  weight_matrix_layer1_type := (
  0 => (-4, 16, -19, -2, -6, 12, -12, 6, 8, 10, 16, -18, -13, 17, -13, 18, -11, 16, -9, -34, -23, 43, 3, -5, -14, 17, 5, -20, 2, -16, -10, 2, -11, -17, 17, 13, 4, -5, -1, 24, 42, 51, 5, 23, 16, -2, -28, -3, -9, 38, 19, 6, 12, -17, 7, -13, 12, 20, 9, -3, 18, -12, 12, 7, -18, 11, -6, 44, 3, 19, -8, -20, -48, -72, -27, -20, 38, 31, 96, 112, 43, -2, 20, 7, 19, -3, -13, 15, 15, -16, 17, 20, -17, 20, 31, 7, 52, 27, -18, -28, -44, 12, 28, 10, 39, 36, 83, 63, 52, 23, 8, 7, 13, -17, 19, 3, 5, -1, 17, -19, 23, 21, 19, 41, 40, 23, -14, -40, 2, -2, -1, 5, 39, 80, 72, 72, 22, 0, 6, -2, 12, -4, -11, -5, -10, -9, 4, -10, -4, -6, -9, 3, 15, 14, 11, -8, -14, 8, 31, 16, 7, 45, 59, 36, -6, 7, -6, 20, -18, -14, -4, 4, -11, 15, -5, -2, -21, -79, -23, 8, 1, 6, -1, -20, -14, 18, 14, 6, 9, 31, 28, 12, -24, 3, -1, 6, 19, -14, 10, 15, 0, 16, -14, 11, -31, -6, -28, -21, -25, -38, -17, -22, 17, -8, 15, 9, 43, 68, 30, -13, -6, -16, 6, -3, 19, 17, -13, 14, 5, 16, -14, 38, 7, 8, 15, -10, -36, -48, -12, -4, 20, 1, 9, 18, 7, 21, 11, -35, -3, -42, -27, -17, -3, 15, -10, -20, -5, 18, 37, 15, 55, 3, -23, -48, -35, -18, -7, 21, 21, 20, 16, 35, 14, -1, -45, -22, -40, -11, -46, -13, -19, -6, -10, -19, 16, 44, 10, 39, 18, -1, -51, -26, -29, -31, -7, 17, 45, 39, 30, 38, 24, -21, -33, -42, -50, -26, -27, 28, 16, -15, 0, -18, -2, 26, -3, 7, -24, -13, -42, -57, -57, -37, -12, 39, 29, 31, 8, 26, -10, -18, -11, -82, -80, -39, -12, 36, 5, 3, 8, -6, 15, 45, 9, 10, -58, -32, -96, -42, -57, -26, 43, 59, 23, 3, 40, 23, -3, 21, -18, -24, -15, -67, 5, 36, -7, 8, -20, -20, 12, -13, -18, -40, -80, -98, -57, -79, -63, 14, 46, 55, 29, 4, 6, 29, -12, 7, -24, 6, -18, -51, -27, -9, 3, 3, 3, 21, 13, -7, -35, -58, -134, -108, -79, -55, -53, 25, 56, 55, 5, 19, 23, -19, -25, -7, -18, -5, -24, -65, -23, -18, 15, -13, -20, -20, 6, -16, -26, -93, -111, -43, -42, -47, -32, 25, 55, 50, 17, 16, 6, 7, -22, -21, -49, -36, -25, -35, -10, 5, 3, -9, -13, -5, -22, -4, -21, -70, -51, -28, 4, -12, 6, 44, 16, 29, 22, 15, 6, 26, -12, -59, -40, -28, -14, -52, 20, -3, -20, -18, -15, 3, -10, -8, -41, -63, -35, -16, -18, -37, 39, 46, 54, 18, 39, 33, 19, -11, -13, -18, -45, 11, -12, -29, -8, -17, -3, 6, -15, 21, 5, -37, -64, -73, -26, 20, 7, 17, 35, 36, 46, 54, 37, 13, 17, 9, 21, -10, -26, 15, -28, -54, -7, 34, -11, 20, 7, -18, -58, -136, -79, -37, -25, 33, -4, 44, 32, 36, 50, 37, 24, 35, 40, 18, -3, -48, -43, -12, -4, -14, -11, 20, -17, -17, 2, 20, -17, -89, -43, -58, 0, -17, 32, 60, 57, 41, 67, 10, -11, -22, -23, -9, -31, -34, -53, -27, -18, -9, -20, 33, 10, 2, -1, -20, 8, -60, 9, -19, 12, 18, 56, 86, 82, 38, 32, 4, 23, -13, 14, -29, -12, -47, -10, -55, -32, 13, 5, 8, -20, 12, 6, 13, -12, 3, 11, 23, 34, 41, 43, 68, 72, 29, 47, 15, -6, 22, 7, -12, -28, -29, -11, -38, -29, -9, 23, 12, -3, -5, -18, 8, -1, 5, 19, 16, 26, 26, 34, 30, 25, 25, 20, 26, -3, 7, 12, -26, -33, -50, -49, -3, -20, -11, -14, -30, -7, -9, 19, 16, -26, 6, 37, 27, 49, 32, 14, 35, 29, 24, 7, 48, -20, -18, -1, -20, -46, -55, -27, -4, 11, 3, -14, 0, 18, -18, -8, -4, 7, 26, 37, 44, 15, 16, 6, 48, 13, 2, 13, 34, 5, -9, -29, -58, -84, -60, -42, -9, 4, 0, 7, 21, 15, -4, -13, 19, 18, 10, 66, 17, 24, -39, -8, -29, 4, -5, 25, -9, -32, -47, -37, -55, -76, -77, -70, -41, -15, -31, -3, -41, 17, -18, 2, -11, -20, 21, 29, 7, 37, -6, -5, 24, 28, 11, 16, 13, -38, -19, 10, -15, -32, -26, -22, 9, -5, -22, -9, -16),
  1 => (-6, -4, 18, -8, 6, 11, -11, -11, -16, 17, 2, -14, -5, 15, 21, 10, -4, 0, -5, -6, 1, 20, 5, 15, 10, 8, -1, -3, -2, 19, 10, -17, -5, -12, -17, -15, 13, -12, 11, -7, -6, 5, 6, 1, 9, -26, -19, 11, -17, -14, 5, 7, -3, 5, -3, 14, 3, 10, -18, 0, 19, -9, 1, 12, 12, -14, 1, 12, -18, -7, 12, -2, 3, 5, -35, -31, -17, -5, -4, -16, -5, -19, -11, 9, 3, -16, 4, -8, 16, 5, 3, 12, -14, 9, 8, -1, -34, 13, -61, -60, -22, -13, -7, -13, -60, -26, -25, -35, -2, -9, 19, -20, 20, 4, -19, 20, 0, -1, 5, 6, 4, -18, -38, -38, -42, 8, -29, -39, -33, -27, 8, 8, 22, -6, -7, -2, 12, -13, -19, -12, -3, -7, 2, -8, -19, -20, 0, 6, -7, 1, -25, -53, -55, -50, -41, -4, 4, -7, 26, 29, 2, 18, -11, -41, 2, 2, -7, 8, -4, 8, 7, -16, 15, -20, 17, 2, -16, -19, -8, -4, -33, -29, -23, -6, -2, 21, 23, -7, 2, -5, -19, -31, -45, 23, 3, 20, 15, 10, -8, -7, 16, 14, -21, -19, 25, 41, 20, -8, 4, 1, -3, -24, -6, 13, 7, -7, 13, 6, -5, 8, -11, 34, -22, -7, -3, 0, -1, -19, -3, -17, -13, -44, 33, -4, 17, 8, 6, 13, 0, 38, -4, -35, -10, -9, -11, 25, 3, -14, 4, 22, -6, -3, 13, -3, -2, -8, -15, 19, -12, -20, 51, 36, 16, 1, 10, 2, 15, 21, 23, -33, 1, -12, -1, -3, 31, -14, 1, 15, 36, 21, -20, -19, 15, 20, -5, 21, -7, -6, -16, 7, 22, 30, 5, 3, -24, -3, -19, -5, 5, -18, -43, -47, 23, -29, -7, -6, 27, 24, -14, 4, 0, -18, 13, 11, -31, -20, -15, -2, 10, 18, -9, -29, -5, -35, -12, -18, -6, 11, 1, -25, -20, -17, -6, -10, 18, -17, -5, -10, 2, -5, -20, -5, -32, 10, 2, -14, 7, 16, -7, 17, -7, -22, -1, 3, -1, 11, -5, -5, 10, 17, -15, -12, -65, -10, 13, -3, -1, -6, -16, -26, -1, 18, 47, 2, -5, -18, 5, -10, 7, -3, -23, 2, 5, 4, 4, 21, 1, 17, 7, -42, -19, -12, 5, 4, 4, 3, 7, -31, 18, 5, 11, 15, -6, 5, -16, -6, -27, 0, -11, -20, -23, -16, -21, 9, 11, 18, 24, -40, 15, 1, -15, 12, 0, 5, -12, -28, -24, -23, 0, -5, -11, 33, -13, -10, -31, -4, -24, -18, 9, -3, 9, 7, 21, 3, 25, -11, 44, 11, -8, -11, -11, 1, -5, -7, -81, -49, -69, -62, -60, -18, -41, -40, -42, -63, -67, -40, -18, 0, 16, 8, 23, 27, 22, 25, 56, 29, -10, -1, -19, 18, 6, -23, -65, -107, -133, -170, -97, -121, -78, -71, -53, -53, -33, -20, 0, 14, 40, 35, 71, 51, 25, -26, 33, 43, 16, -11, 1, -8, -1, -12, -94, -77, -99, -139, -99, -79, -62, -15, 20, 38, 8, 47, 59, 44, 23, 17, 14, 44, 0, -8, 3, 1, 12, -13, -5, 12, -7, 1, -22, -18, -13, -18, -7, 33, 31, 48, 38, 52, 42, 25, 32, 24, 18, 25, 7, 15, 28, 15, 7, -42, -6, -7, -1, 15, -25, 28, 10, 24, 43, 34, 88, 47, 64, 57, 46, 33, 21, 40, 53, 18, 8, 26, -9, 25, -5, -3, 6, -2, -1, 17, -15, 20, 17, 32, 11, 45, 41, 66, 39, 24, 42, 33, 21, 57, 43, 68, 34, 18, -14, 6, 27, -17, -5, -5, 11, 18, -14, 6, 1, 11, 10, 27, 41, 57, 56, 61, 52, 49, 63, 25, 32, 58, 26, 37, 10, -3, -23, -41, -21, -66, -51, -36, 33, 57, 4, -13, -3, 14, 34, 39, 16, 22, 71, 27, 25, 40, 26, 65, -1, -2, 21, -9, -9, -51, -46, -26, -26, -29, -66, 15, 53, -3, -1, 6, 11, -15, 45, 25, 59, 8, 40, 28, -8, 4, 5, 1, -8, 0, -46, -43, -23, -57, -23, -32, 5, -9, -14, -2, 8, -7, 18, 1, 19, 17, 8, 1, -13, -10, 12, 0, -37, -26, -34, -35, -70, -70, -51, -10, -11, -36, -67, -45, -46, -12, 53, 3, 0, 7, 6, 17, 10, 4, 0, -32, -45, 17, 4, -6, -7, 19, -4, -49, -54, -50, -36, -66, 2, -30, -14, -24, -50, -45, -18, -6, -8, 2, -1, -11, 5, -12, -17, 13, -15, -23, 23, 31, 7, 5, 28, 55, 17, 37, 14, -37, -31, -24, -24, -29, -33, -9, -24, -5, 43, 7),
  2 => (-20, -11, -11, -7, 15, -17, -11, 6, 9, 6, -1, -20, 14, 20, -4, -24, -57, -11, -9, -4, -13, 26, -18, -13, -15, 19, -1, 8, -13, 2, -14, -3, 6, 12, 5, 7, 12, 7, -10, 23, -31, -2, 10, 19, 9, -29, -38, -37, -18, 10, 25, -1, 32, 18, 1, -19, -9, -8, 1, -7, -13, 14, 11, 18, -1, 20, 3, -26, 24, -33, -31, -19, 18, 79, 3, 42, 21, 38, 32, 58, 20, 25, -7, -12, 19, -16, 3, 17, -13, -3, 20, -4, -1, -12, 3, -7, 4, -16, 2, -24, -24, 4, 3, 44, 39, 50, 25, 2, 9, -9, -4, 12, -7, 6, 0, -11, 4, -6, 5, -15, 47, 80, 49, 49, 27, 10, 5, -8, 20, 35, 35, 14, 11, -14, -2, -41, -12, -17, 6, -2, 14, 16, 15, -4, 10, -14, -37, 6, 33, 31, 24, 21, 13, 26, 42, 10, 50, 23, -8, -57, -54, -35, -47, -77, -34, 16, -13, -6, 9, -16, -16, -9, 10, 13, -10, -41, 34, -17, -30, -16, -46, -22, -38, -48, -54, -89, -111, -134, -149, -110, -69, -78, -26, 2, 22, 2, -18, 5, -1, 6, 9, 5, -28, -37, -26, -19, -60, -4, -24, -17, -14, -24, -21, -17, -50, -68, -33, -39, -38, -50, -2, -13, -35, -28, -9, 16, -2, -20, 5, -3, -41, -19, -16, 4, 59, 36, 13, -8, 6, 15, 19, 10, 15, 29, 27, 37, 69, 31, 21, -14, -40, -17, 3, 2, -5, 11, 2, 15, -54, -21, 39, 20, 42, 70, 34, 18, 8, 9, 10, 17, 23, 26, 28, 27, 21, 76, 38, 18, -5, -27, 14, -11, -15, 13, -15, -22, -46, -24, 3, 18, 20, 25, 8, 10, 42, 39, 37, 64, 49, 57, 39, 47, 45, 33, 43, 39, 35, -14, -19, 19, 2, -3, 11, -14, -44, -22, -16, -54, -65, -65, -67, -82, -42, -17, -10, -19, -27, 7, -1, 29, -8, 12, 35, 29, 10, 7, -8, -15, 14, 1, -18, -27, -9, 7, -32, -43, -69, -48, -88, -82, -58, -65, -81, -94, -82, -66, -52, -55, -46, -18, -20, -6, 21, 28, -6, -10, 17, 15, -4, -19, 0, 7, -18, -35, -17, -7, 11, -16, -20, -32, -46, -35, -80, -53, -34, -45, -28, -49, -62, -26, -29, 4, -13, 14, -6, 8, -17, -17, -18, 11, 28, 35, 60, 37, 58, 33, 34, 17, 14, 35, 38, -15, -23, -36, -29, -34, -85, -61, -15, -2, -17, -17, 6, 7, 9, -17, -30, -14, 29, 35, 28, 24, 45, 28, 22, -5, 4, 20, 13, 13, 24, 2, -6, -53, -68, -72, -49, 0, 13, -10, -4, 0, -23, -9, -20, -8, 26, 25, -9, -4, -13, 5, 17, 19, 13, 11, 6, -6, 21, 6, -8, -22, -17, -50, -42, -34, 13, 9, -9, 0, -10, 31, 17, 33, 25, 27, -9, -8, 6, -28, 9, -17, 28, 31, 42, 7, 0, -12, 8, 3, 12, -5, -5, -6, -2, 12, 3, -7, -37, -19, -12, 12, -27, -35, -49, -18, -29, -52, -15, -26, -51, 0, 9, -4, -35, -17, 4, 18, 15, 12, -6, -8, 19, 12, -5, -5, -38, -77, -24, -14, -14, -2, -11, 0, 17, 25, -2, -18, -40, -46, -15, -19, -7, -20, -26, -8, 31, 17, 20, -9, -6, 10, 9, 13, 1, -47, -33, -30, -25, 14, 48, 57, 13, 54, 62, 53, 23, 8, 14, 11, 24, -6, 1, -27, 27, 13, 34, -26, 8, -4, 5, 6, 0, -38, -28, -31, -18, -5, 4, 19, 20, -13, 7, 2, -14, 22, 3, 25, 18, 6, -12, -23, -14, -26, 18, 6, 19, -7, 2, 16, 8, -4, 8, -26, -29, -4, -29, 2, -14, -4, 0, -14, -21, -9, -5, 1, -16, -14, -14, -4, -28, -17, 0, -38, -16, -12, -6, 4, 10, 9, 14, 16, 0, 13, 28, -4, 0, 20, 11, 25, -27, -16, 12, -8, 3, -17, 8, -6, -5, 4, 13, -25, -18, -15, 5, 11, -31, -11, 3, -18, -28, -10, -12, -9, 4, -29, -13, 14, 14, -8, -16, -27, 0, -39, -32, 30, 2, 6, 23, -26, -1, -13, -16, -5, 13, 22, 2, -25, -26, -32, -28, 28, -2, 8, -33, -44, -1, -35, -11, -9, 4, 7, 28, 21, 18, 31, 12, -5, -12, 15, -2, 15, 11, -1, -21, -8, -12, -39, 1, -12, -38, -27, -48, -23, -47, -35, 16, -29, -40, -9, 11, -11, 8, 7, 8, -10, -16, 20, -3, 17, -15, -8, -7, 2, -7, -29, -27, -29, -16, -20, -20, 5, 18, -17, 2, -11, -41, -40, -39, -43, -11, 22, -4, -9),
  3 => (-7, 3, 15, -19, 20, 9, 3, 3, 17, 4, -13, 21, -4, 18, 40, -4, -19, -4, -35, -6, -36, 39, -3, 20, -7, 15, -7, -1, -4, 5, 18, -2, -15, -4, 5, 18, 0, -5, 13, -5, -22, -23, 19, 2, 21, 50, 24, 40, 42, 8, 28, -21, 0, -6, 3, 16, 4, 2, -15, -6, -3, -21, 0, -14, -15, -9, 26, 26, -3, 2, -25, 3, 8, 6, 1, 31, 54, 51, 34, -10, -9, 17, -13, 4, -17, 2, 4, 13, -20, 12, -13, 18, 10, 23, -15, -30, -27, 18, -17, 2, 30, 2, 27, 35, -2, -13, 3, 41, 5, 1, 6, -21, -13, -12, -19, 10, 6, 5, 20, 26, 6, 8, -7, 4, -16, -10, -11, -33, -4, 17, -6, 12, 0, 5, 28, 28, 13, -10, -5, -3, -6, 10, -5, -2, 0, -7, 32, 29, 58, -20, -7, -5, 6, -29, -13, 15, 17, 34, 39, 3, 16, 28, 7, 46, 18, -13, 6, -19, 4, -5, -9, 9, 5, -13, 12, 67, 19, -5, 9, 30, 48, 42, 10, -7, 33, 52, -11, 1, 4, 37, 47, 39, 55, 35, -4, -8, 10, 1, 15, -3, 0, 9, 15, 44, 58, 65, 42, 67, 64, 64, 15, 15, 38, 43, 26, 19, 44, 37, 49, 43, 37, 34, 65, 18, -12, -7, -8, -11, -12, 5, 25, 62, 91, 72, 72, 104, 81, 24, 33, 34, 43, 52, 50, 16, 31, 70, 59, 60, 75, 77, 84, 45, -14, 4, -3, 19, 10, -8, 26, 82, 75, 106, 84, 86, 54, 65, 70, 51, 32, 36, 35, 36, 41, 21, 19, 20, 58, 86, 49, 21, 17, 20, 4, -5, 19, 48, 60, 61, 71, 59, 61, 81, 83, 58, 56, 27, 66, 50, 3, 15, 47, 19, 49, 33, 45, 92, 63, 41, -8, 15, -9, 8, -14, 34, 73, 32, 77, 74, 66, 75, 82, 75, 46, 62, 58, 30, 22, 32, 17, 18, 33, 35, 36, 59, 82, 50, -17, -5, 2, 16, 24, -4, -6, 5, 60, 27, 20, 45, 40, 35, 32, 7, 39, 10, -5, 23, 2, 19, 54, 4, 3, 59, 38, 42, -18, 10, -3, 9, 30, -12, -16, 21, 32, 31, 34, 41, 35, 24, 14, -4, -3, 12, 28, 9, 29, 57, 52, 14, -37, 38, 37, 20, -8, 3, -19, 21, -8, -5, -15, -11, -12, 21, 31, 11, 35, 10, 23, 12, 32, 39, 58, 63, 5, 39, 51, -11, -10, 7, 36, -1, 10, -2, 9, -18, 15, -17, -18, -52, -47, -34, -22, 7, 11, 10, 14, 18, 59, 40, 66, 23, 0, -8, 7, -4, -34, 23, 8, -4, 6, -12, -10, -2, 23, 3, -35, -59, -35, -37, -13, -8, -4, 21, 42, 16, 38, 29, 37, 14, 5, -16, -15, 4, -1, -8, -3, -6, 17, 11, -7, 2, -20, -25, -43, -51, 4, -42, -40, -16, 9, 2, 39, 59, 20, 19, 9, -2, 3, -18, 3, -30, 7, 11, -19, -3, -12, -5, -6, 9, -17, 5, -15, -18, 7, 13, -26, -17, 34, 31, 16, 46, 5, 18, 9, -17, -9, -10, -13, -33, 11, -2, 10, 26, 17, 5, -8, 17, -25, -6, 15, -7, -2, -17, 18, 25, 21, 40, -25, 19, 12, -27, -5, -11, 8, 17, 0, -44, -44, 7, 22, 12, 3, 7, 18, -12, 5, -31, -25, -22, -44, -10, 12, -36, -20, 1, -6, 10, 5, -7, -11, 0, 18, 35, 33, -1, -33, -1, -13, -27, -14, -5, 2, -13, -13, -21, -32, -36, -22, -45, -4, -40, -16, -28, -18, -17, 10, -6, 16, 32, 3, 9, 16, 0, -17, -4, -15, -22, -2, 9, -6, 21, -27, 13, -42, -34, -15, -59, -8, -53, -34, -13, -2, 22, -3, 7, -11, 9, 2, 29, 7, -15, -1, -6, -29, -16, 14, -15, 17, -16, -39, -22, -5, -3, -15, 5, -19, -39, -13, 21, 30, 27, 49, 34, 10, -35, -15, -10, -2, 10, 7, -3, -49, -9, -18, -14, -20, 4, 6, -11, -9, 6, 9, 45, 36, 3, -16, 12, 5, 52, 13, 20, -18, -15, -20, -23, -2, -11, 15, 5, -24, -74, -19, 18, -5, -18, 35, 44, 68, 23, 16, 43, -11, -13, 6, 18, 32, 17, -5, 34, -13, -8, -1, -29, -8, 30, 16, 20, -23, -51, 0, 9, 18, -9, 18, 52, 49, 37, 28, 44, 38, 9, 43, 35, 56, 24, 38, 35, -15, -28, -2, 23, 54, 35, 37, 18, -23, -22, 14, 7, -8, 12, -20, 35, 30, 83, 102, 81, 53, 68, 37, 42, 86, 35, 37, 58, 8, -30, 41, 45, 42, 50, 12, 4, -11, -32),
  4 => (21, 14, 4, 1, -4, -18, -15, 16, -5, 19, -3, -14, -17, -21, -4, 6, 6, -29, 8, 24, 28, -28, 10, -16, -16, -1, 13, -5, -11, 7, 21, 4, 12, -1, 13, 5, 8, 14, 22, -4, -17, -5, -9, 4, -10, 8, 26, 14, 36, 46, -32, -10, -10, 8, 17, -13, 9, 20, -6, 9, -13, -12, 18, 11, -2, 11, 28, 14, 29, 21, -10, 19, -17, -7, 31, 28, -11, -5, -46, -24, -16, 19, -15, -5, -19, 10, -20, -18, -11, -17, 14, 16, -12, -12, -20, -32, -47, -33, 13, 13, 19, 26, 28, 17, 18, 28, -20, -12, 26, 17, 3, 16, -12, 15, 12, 20, -7, -19, -10, -3, -23, -98, -86, -116, -53, -24, 0, 4, 5, 52, 64, 24, 38, -6, 0, -10, -9, 11, -20, -10, 3, -12, -13, -13, 11, 19, -38, -11, -49, -61, -92, -110, -46, 8, 10, 3, 5, 46, 20, 44, 18, 11, 1, -17, -38, 21, 19, 0, 7, 18, -16, -13, -8, -20, -48, 6, -9, -74, -97, -56, -14, 8, 26, 36, 31, -6, 45, 20, 35, 31, 3, 2, -14, -16, 20, -12, 19, -10, 8, 19, 8, -17, -25, -1, -5, -103, -98, -32, 15, 51, 20, -29, -9, 15, 17, 4, 8, 7, -6, -23, -4, 6, 7, 20, 2, -6, 18, 8, 19, -10, 4, 28, -2, -75, -49, -8, 46, 29, 31, 0, -8, 0, 28, 25, -5, -5, 1, -34, -18, 5, 35, -1, -18, -2, 2, -19, 0, -15, 68, 56, 5, -43, -27, 43, 39, 37, 59, 9, -11, -30, -11, 14, 19, 9, 32, 31, -40, -28, -6, 2, -16, -20, 2, 5, -12, -13, 54, 64, 6, -30, -6, 60, 52, 66, 39, -3, -15, -64, -3, -6, 11, -5, -25, 33, -40, -54, -61, -11, -13, 5, 7, 0, 8, 31, 82, 37, 6, -26, 39, 64, 64, 23, 12, -44, -53, -42, 11, -13, -40, -55, -10, 10, -30, -74, -45, 3, 11, -14, 20, 5, 14, 27, 32, 6, -15, -9, 33, 80, 71, 37, 46, -43, -48, -50, 16, -24, -31, -30, 3, -9, -55, -53, -41, 18, 3, -12, -6, -14, -5, 4, 10, 13, -48, -5, 32, 32, 72, 67, 6, -41, -49, -31, 15, -5, -2, 7, -12, 6, -30, -81, -13, -11, 15, 10, 9, -19, 0, 37, 13, -50, -79, -21, 29, 43, 20, 7, -1, -51, -67, -15, 5, 36, 2, -13, 15, 13, -40, -48, -13, -1, -8, 12, -9, -16, 1, 2, -17, -44, -85, -31, 4, 27, 34, 15, -31, -55, -36, -35, 3, 29, 17, -4, 18, -4, -46, -28, -39, -38, -7, -4, 16, 6, 31, 10, -17, -45, -74, -30, 35, 15, 32, 25, -32, -53, -62, -53, 8, 11, 8, 25, 19, 7, -28, -31, -49, -13, -9, 0, -7, 18, -18, -27, -69, -85, -86, 4, 33, 24, -4, 10, -24, -76, -54, -30, -10, 0, 23, 19, 15, 21, -40, -73, -25, -39, -2, 16, 13, 12, -44, -48, -81, -119, -88, -52, 17, 8, -21, 10, -10, -56, -5, -19, -19, 29, -3, 4, 17, 0, -24, -69, -12, -2, 3, -11, 3, -14, -23, -38, -112, -120, -136, -37, 30, -23, 3, 19, 0, -21, -46, -27, -26, 22, -15, 12, 35, 16, -94, -42, -25, -5, 17, 19, 20, -11, -44, -58, -85, -118, -128, 4, 30, -2, 24, 19, -25, -20, 25, 21, 13, 10, -33, -17, 20, -43, -84, -46, 11, -21, 19, 17, 15, 18, -28, -58, -90, -104, -122, -31, 41, 37, 16, 34, -16, 4, 8, -27, -41, -11, 13, -11, 53, -18, -72, -68, 2, -2, 8, -1, 7, -5, -5, -42, -42, -102, -101, -64, 27, 36, 45, 29, 18, -25, 10, -23, 2, 6, 40, 18, 31, -45, -66, -21, -42, 11, 18, 4, -2, 9, -28, -55, -53, -50, -74, -70, 1, 47, 19, 31, 15, -13, -3, -13, 29, 24, -2, 23, 1, -70, -71, -46, 1, -8, -17, 1, 0, -14, 5, -43, -47, -28, -49, -61, 2, 6, -5, -5, -9, -15, -4, 36, 22, 18, -7, 18, -39, -66, -8, 13, 10, -1, 5, 1, 6, -14, -22, -19, 1, -6, -14, -17, -3, -17, -16, 0, -27, 5, 32, 18, 8, 24, 20, -22, -49, -65, -33, -19, -25, -35, -2, 6, -19, 16, -16, -1, -27, 8, 7, 0, 25, -36, -7, 1, -37, -28, 11, 18, -15, -29, -29, -32, -49, -46, -100, -40, -44, 8, -13, -1, 18, 19, 9, 15, 5, 7, -15, 0, 2, -25, -30, -2, 9, 8, 27, 33, 33, 23, -23, 3, 13, -23, -33, -21, -24, -22),
  5 => (-10, -14, 20, -15, -15, 0, -16, -6, 14, -13, -20, -17, 20, -13, 8, -13, 23, -4, -34, 9, 52, 28, 6, -17, 16, -7, -8, 19, -7, 3, -12, -9, -1, 19, 4, 15, 14, 12, 34, 2, 12, -10, 62, 70, 66, 55, 46, 17, 94, 75, 48, -34, -9, 5, 3, 21, -17, 8, 15, 8, -11, -12, -7, -19, 8, -1, -21, 26, 30, 46, 42, 47, 54, 65, 9, 9, 41, 43, -5, -69, -21, 14, 9, -18, 10, -17, 10, 14, -4, -6, -17, -14, -16, -33, 5, 72, 64, 47, 0, 44, 36, -17, -9, -2, -17, -6, 37, -10, 13, 27, 17, 13, 17, 4, -17, 1, -20, 17, 18, -11, -10, 10, 41, -13, -24, -34, -26, 16, 15, -23, -19, -22, -24, 0, 38, 7, 35, 22, -1, 10, -13, -4, -4, 4, -11, 4, -34, -41, -41, -38, -32, -57, -22, -10, 31, 27, 0, 9, 40, -7, -3, 46, -2, 50, 30, 10, -7, -11, -10, 19, -5, 19, -19, -9, -68, -48, -42, -6, -4, 18, 29, 34, 49, 53, -1, 22, 48, 36, 61, 67, 57, 29, 43, 7, 19, -10, 0, 3, -20, -5, 19, -7, -46, -8, -13, 44, 64, 18, 1, 35, 24, 13, -27, -6, 33, 17, 47, 62, 39, 26, 13, -2, 44, -5, 7, 15, -20, 5, 18, 0, 11, 52, 48, 78, 22, -14, 4, 32, 38, 12, 6, 6, 38, 16, 27, 37, 38, 10, 3, 51, 64, 42, 12, -7, 11, 4, 17, 13, 44, 45, 47, 85, 33, -3, 33, 11, 24, 39, 26, 54, 17, -1, 17, 26, 42, -7, -16, 31, 69, 51, 11, -18, -7, 16, -6, 0, 55, 71, 58, 60, 38, 50, 46, 20, 33, 36, 39, 38, 5, -38, 3, 26, 21, -15, -5, 32, 47, 60, -2, 11, -6, -2, -1, -1, 104, 96, 85, 79, 90, 85, 80, 47, 43, 59, 62, 54, -3, -2, 19, 63, 48, -12, 8, -28, 8, 62, -10, -13, -2, 9, -21, -6, 85, 54, 89, 97, 93, 93, 69, 60, 74, 95, 75, 50, 53, 40, 13, 48, 32, 28, 10, 1, 7, 49, -10, 8, -20, -11, -27, -7, 16, 63, 68, 57, 44, 56, 26, 40, 50, 37, 47, 25, 36, 12, 65, 85, 47, 45, 10, -34, 2, 38, 3, 16, 5, -16, -22, 28, 41, 37, 6, -8, 23, 5, -36, -31, 41, 43, 28, 46, 37, 45, 33, 22, 36, 8, 53, -16, -15, 7, -7, 17, -13, 4, -6, 41, 70, 10, 18, -31, -2, -4, -33, -1, 6, 40, -4, 41, 58, 16, 38, -11, 25, 21, 2, 25, -40, -38, 15, 17, 11, 17, 18, 10, 12, -17, 12, -3, 7, 26, 37, 15, 59, 19, 4, 44, 49, 19, 46, 5, -13, -6, 7, 12, -17, -35, 11, -11, -9, 4, -14, -23, 3, -42, -34, -24, -5, -7, 7, 22, 51, 20, 15, 0, -15, -3, 4, 12, 2, -16, 25, 17, 11, -6, 16, 14, -4, -19, 16, -16, 14, -29, -37, -29, 7, 15, 41, 21, 19, 41, 27, 36, 19, -32, -8, -1, -13, -28, 9, 47, 48, -21, -7, -3, 20, -2, 20, 5, 11, -27, 6, -20, 2, -5, -10, 5, -9, 11, 4, 7, 3, -39, 13, 13, 4, -12, 4, 19, 9, -7, 9, 2, 11, 0, -39, -35, -63, -65, -49, -15, -8, -31, -12, -18, -28, 7, 16, -10, -8, -30, 29, -4, 10, -15, -21, 17, 6, -9, -9, -18, 5, -5, -17, -2, -34, -49, -39, -19, 0, 3, 0, -13, -26, -4, 5, -19, -13, -17, 5, 14, 7, -13, 25, 38, -2, -6, -11, 12, -8, -15, -16, -10, -26, -32, -50, -47, -5, -54, -25, -14, -38, -20, 5, -10, -1, -13, 0, 19, 7, 22, 20, -5, -34, -69, 3, -3, 1, 1, -31, -60, -54, -36, -30, -31, -16, -3, -6, -19, -11, -4, -4, -3, 16, -13, 8, -3, 0, 33, 43, -33, -30, 7, 18, -3, 20, 12, -23, -38, -31, -39, -26, 8, 32, 22, 29, -12, -13, -14, -21, -27, 8, 5, -26, -28, 3, 14, 40, 2, -7, 2, 16, 6, -5, 17, 43, -21, 11, -13, -21, 29, 43, 39, 19, 18, 9, 15, -12, 7, -15, -7, 12, 18, 6, 19, 47, 14, -6, -10, 13, -1, 19, 6, 20, 9, 10, 17, -10, 35, 69, 21, 56, 81, 60, 56, -19, 18, 32, 0, 8, 1, -29, -2, -4, 33, -19, -15, -16, 0, 0, 7, -16, 12, 21, 47, 36, 31, 72, 72, 56, 60, 53, 36, 62, 63, 0, -17, -20, -3, -5, -3, 14, 21, -12, 9),
  6 => (-12, 10, 21, -14, -1, -8, -4, -1, 12, 1, -19, 10, 7, -10, 20, 4, 9, 41, -8, -38, -10, -1, -10, -5, 12, 14, -19, -1, 9, 2, -15, 13, 5, 11, -5, 19, -8, -7, 7, 33, 46, 2, 5, 29, 61, 62, 22, 7, 12, 17, 29, 36, 27, -15, -13, 19, -20, -3, -9, 11, 15, 15, 12, -16, -5, 14, 0, 15, 32, 74, 105, 76, 39, 69, 57, 20, 31, -14, 7, 38, 36, 13, -19, 19, -21, 8, -14, -16, -15, -11, 12, -14, -5, 35, 10, 30, 38, 43, 46, 14, 34, 24, 21, -19, -7, -24, -2, 12, -12, 10, -4, -15, -3, -10, 2, -10, -11, 8, 16, -39, -23, -95, -38, 11, 11, 53, 68, 38, 24, -19, 9, -9, -5, -14, 33, 10, 15, -25, 16, 16, -9, -7, 10, -5, -6, -20, -19, -51, -82, -17, -5, -2, 22, 31, 25, 23, 32, 20, 3, -1, 5, 30, 33, -31, -46, -35, -11, -4, 3, 4, 16, 1, -4, 2, -58, -16, -50, -25, 10, -42, 10, 10, -3, 5, 48, 40, 22, 3, -3, 4, 26, -12, -41, -45, -22, -16, -8, 3, -8, -14, 20, 2, -19, -6, -37, -3, -52, -44, -1, 6, 54, 63, 45, 31, 37, -19, -9, 4, 20, 0, -15, -6, -32, -2, -17, 11, -5, 1, 10, -3, -18, 26, -23, -24, -8, -15, 4, 40, 63, 41, 20, 35, 14, -35, -47, -44, -38, -26, -24, 24, -24, 10, -17, 16, -4, -2, -16, 8, 42, -2, -46, -17, -16, -2, 50, 57, 93, 54, 3, -16, 14, -5, -5, -3, -11, 7, -37, -40, -37, 4, -3, 19, 1, -3, 1, -43, 33, -10, 13, 18, 34, 23, 17, -10, 25, 12, 22, -13, 28, 11, -4, 32, 24, 26, -12, 3, -14, 2, -14, 9, 0, -17, -15, -66, 26, 18, 21, 50, 56, 55, 24, 16, 39, 13, -2, -19, 28, 16, 9, 13, 15, 24, -7, 18, 3, -40, -19, 16, 5, -5, -16, -23, 84, 84, 75, 77, 62, 63, 14, 33, 45, 39, 29, 12, 37, 28, -1, -26, -9, 13, 9, 20, 13, -11, 19, 21, 9, 14, 23, 8, 107, 127, 97, 58, 86, 69, 15, 35, 70, 60, 26, 39, 43, 51, -4, 4, -6, -7, 32, 35, 5, -48, -14, 20, 0, -9, -36, 6, 92, 95, 71, 70, 55, 41, 13, 41, 29, 34, 43, 25, 1, 24, 43, 25, 45, 52, 67, 95, 45, 5, -7, -7, 7, 19, -33, -13, 58, 28, 4, 45, 21, 10, 0, 21, -16, -2, 13, 0, -5, 2, 30, 22, 70, 80, 93, 98, 49, -18, 4, -4, -18, 20, -33, 19, 33, 21, 0, 16, 14, 1, 8, -6, -17, -18, 3, 7, 22, -9, -33, -1, 19, 58, 110, 96, 59, -22, 18, -4, 8, 10, 1, 31, 51, 12, 30, 26, 4, -28, 8, -7, 11, 1, -15, -16, -5, 17, 56, 5, 28, 102, 71, 92, 88, 43, -14, 15, 8, -2, -11, 16, 21, -22, 5, 5, 36, -2, 8, 18, 21, 10, 9, 22, 13, 25, 59, 53, 48, 73, 48, 56, 74, 24, -3, 3, -14, -20, -11, 11, -9, -19, -34, -28, -10, 44, -5, 11, 8, 31, 29, 20, 7, 12, 36, 18, 44, 52, 27, 49, 37, 1, 15, 17, -10, 2, 5, 24, -24, -14, -20, -32, -13, 6, 27, 36, 25, 46, 57, 56, 69, 66, 72, 33, 23, 50, 0, 34, 12, -19, 5, 9, -2, 7, -20, -27, 38, -24, -14, -8, 49, 36, 33, 49, 62, 43, 28, 63, 38, 84, 70, -15, 21, 28, 10, 5, -3, -3, -2, 15, 17, 1, -42, 15, 2, 33, 51, 18, 33, 19, 27, -8, 1, 21, 12, 18, -5, 31, 38, -23, -4, -14, 10, -13, -37, -44, 9, -6, -7, 8, 2, 11, 10, 25, 20, 32, 4, 29, 21, 3, -45, -25, -3, -18, -9, 0, 2, -17, 20, 14, -6, -15, -46, -41, -10, 0, -2, 7, 2, 17, -18, 27, 5, -18, 10, 3, -21, -19, -15, -32, -16, -24, -8, -6, -23, -11, -19, 2, 11, 22, 9, -13, 1, -3, 19, 20, -5, -13, -5, -8, -28, -37, -20, 0, 2, -19, -18, 9, 23, 23, 3, 10, -19, -7, 2, 5, 15, 53, 26, -15, -7, 14, 5, 19, 3, 49, -27, -30, -4, 2, -8, -25, -18, -17, 2, -34, 28, 6, 41, 11, 6, 17, 13, -9, 17, 1, -25, -11, 10, 9, -19, 12, -19, 44, 29, 19, 38, 25, 19, 13, 43, 38, 43, 25, 36, 61, 71, 7, 40, 3, -2, 14, 24, -4, -7, -52),
  7 => (2, -14, -1, -15, 15, -19, 10, -3, 13, 3, 20, -2, 0, -10, 5, 6, -18, -59, -54, -18, -36, -38, -20, 5, -6, -3, -1, 14, 16, 18, 4, 7, -12, -7, -18, -2, -6, -11, 60, 37, 34, 31, 24, 21, 10, 6, -75, -56, -68, -34, -7, 59, 44, -4, 16, 13, 5, -19, -8, -4, -16, 17, -9, -7, 16, 28, 21, 9, 19, -12, -36, -20, 12, 54, 5, 21, 59, 30, 49, 97, 71, 16, 15, 3, 12, -14, 20, -3, 10, -20, 3, -20, 2, 37, 54, -5, -29, -25, -6, -30, 21, 56, 36, 39, 45, 49, 38, 80, 28, 54, 8, -16, -20, -14, -7, -2, -6, -21, -10, 26, 32, 77, 17, 28, 33, 6, 0, 20, 30, 47, 13, -18, -52, -42, -33, -17, 8, 9, 15, -10, 5, 9, -14, 15, 4, 15, -41, -15, 12, 12, 5, -33, -12, 4, 7, -2, -11, -28, -60, -58, -56, -61, -53, -60, -20, 8, -5, 15, 6, -4, 16, 19, -15, 8, -23, -4, 14, 1, 17, -44, -16, -24, 31, -5, -33, -61, -62, -92, -81, -113, -87, -66, -33, -3, 10, 8, -9, -20, 9, -11, 20, 10, -44, -15, -18, 11, 24, -30, -34, -39, -31, -18, -47, -38, -5, -43, -84, -72, -49, -68, 10, -3, 14, 12, -11, -12, 18, -17, 14, -3, -27, -21, -10, 38, 35, -24, -56, -31, -54, -14, -38, -61, -51, -68, -26, -14, 21, 8, 29, -28, 0, 37, -6, -13, -8, -2, -16, 2, -59, -14, -24, 12, -12, -7, -16, -37, -37, 4, -49, -13, -11, -2, 18, 44, 62, 63, 38, 16, -5, 36, 6, -5, 17, -7, 0, -20, -66, -49, -19, 10, -4, 9, 30, 5, 6, 12, 9, 62, 30, 63, 42, 57, 52, 33, -4, -1, -12, 30, 5, 3, 8, 8, 18, -54, -79, -64, -22, -13, -6, 38, 85, 49, 29, 28, 39, 72, 71, 67, 36, 65, 40, 30, -13, -50, 4, 2, -16, -14, -8, 7, 28, 53, -45, -36, -11, 39, 28, 62, 60, 26, -16, -2, 28, 56, 60, 45, 53, 8, 33, 39, -1, -73, -49, 20, 5, -5, 6, -14, 8, 12, 16, 12, 37, 77, 83, 74, 33, 11, -4, -17, 5, 15, -6, 26, 60, 23, 37, 9, 35, -21, -1, 29, -3, -16, 12, 0, 18, 31, -28, -5, 3, 49, 20, 49, 38, -8, -33, 22, -11, -1, 12, 14, 57, 18, -14, -37, -19, -10, -10, 28, 11, -2, -10, -7, -6, -18, -52, 22, 9, 37, 25, 49, 39, -33, -48, -24, 12, 5, -13, 15, 33, -1, -62, -45, -40, -64, 1, -11, -15, -10, 6, -16, -3, -7, -19, -13, 10, 6, 43, 43, 28, -40, -61, -9, -31, -1, 5, 4, -1, 4, -71, -60, -52, -54, 7, 24, 13, -1, 10, -3, 13, -54, -39, -24, -16, 21, 73, 34, 11, -64, -64, -33, -19, 4, -3, -8, 9, 21, 1, -18, -25, -39, 37, 9, 3, 3, -19, -19, 10, -8, -37, -19, 34, 20, 40, 28, -7, -48, -28, -2, -11, 12, -10, -28, -11, 13, -2, 3, 16, -22, -23, 12, 9, 14, 7, 9, 25, 4, -20, -16, -6, -5, 40, 42, -9, -57, -31, -19, -21, -1, -15, -61, -33, 9, -2, -26, -4, 8, 3, 17, 1, 8, -7, 9, 7, -13, 7, -15, -21, 14, 29, 21, 12, -33, -15, -49, -43, -23, -49, -77, -51, -33, -17, -17, -1, 4, -23, 46, 16, -16, -19, -12, 26, 29, 17, -3, -20, -5, 48, 54, 31, 41, 9, -27, -43, -37, -46, -81, -41, -8, -49, -80, -13, 28, -17, 39, -9, 9, -12, -13, -5, -43, 7, 6, -15, -35, 21, 58, 10, 17, 36, 16, -10, -2, 10, -49, -3, -50, -32, -70, -41, -11, -13, 32, -3, 13, 14, -16, -15, -46, -30, 6, -29, -13, 13, 30, 11, 27, 6, -7, -36, -17, -10, -33, -25, -7, -30, -11, 2, 4, 20, 70, -10, 20, 1, 16, 11, -70, -17, -18, -23, 16, 25, 31, 9, 22, 36, 2, -6, -34, -3, -9, -49, -1, 13, -19, 1, -2, -3, 58, -20, 15, -14, -12, -37, -57, -18, 1, -22, -16, 17, 39, 1, 6, 39, 35, -2, -14, -19, -19, -6, -22, 25, 0, -12, -12, 48, 42, -13, 21, 3, -1, -19, -27, -28, -26, 2, -9, 6, -19, -13, 10, 8, 13, 2, -7, -17, -35, -55, -28, -34, 0, -14, 11, 82, 56, 11, 6, -11, 8, -8, -11, 15, -37, 13, 5, -18, -26, 15, -7, -15, -55, -42, -42, -33, -37, -27, 4, -23, -31, -27, -3, 29, 64),
  8 => (-1, -18, -20, -15, 19, 1, 2, 7, -5, 10, -8, 17, -2, 12, 4, 7, 12, 6, -12, 0, 16, -5, -5, 20, 16, -6, -19, -17, 10, -7, -5, 15, -5, -2, -4, -1, 13, 4, -6, -18, -26, -14, -45, -31, -31, -30, -53, -53, -29, 4, -24, 4, -4, 20, 11, 12, -14, 6, -19, 16, 1, 4, 1, 6, -9, 11, 18, -15, -12, -24, -8, -36, -52, -16, 7, -24, -23, -27, 10, -15, 5, 2, -19, -18, 20, 0, -6, -13, 3, -13, -4, -15, -2, -15, -28, -36, -9, -35, -48, -36, -49, 4, -22, -17, -33, -53, -34, -12, 9, 23, 9, -13, 2, -16, 5, -11, -1, 15, 6, 0, 3, -24, -7, 37, -33, 2, -36, -24, -38, -8, 16, -19, -13, -19, -52, -8, 2, -7, -8, -5, 3, -13, -8, -9, -8, -6, 9, -9, -6, -5, -28, -7, -13, -11, -32, -5, -13, 12, 32, 4, -3, -18, -42, 7, 15, -22, -2, -2, -8, -15, 14, 4, 4, 0, 18, -24, -42, -45, -34, -35, -35, -13, -15, 12, 21, 42, 12, 11, 0, -27, 41, 13, 17, -13, -1, -8, -16, 5, -9, 5, 18, 6, 6, -43, -60, -29, -62, -35, 27, 15, 3, -1, -11, 11, 4, 4, 1, -8, -20, -3, -35, -9, 15, 10, -15, -20, 13, -15, -2, 7, -29, -31, -77, -54, -49, -11, -26, -18, -16, -24, -19, 34, 15, 18, -12, 4, -26, -30, -38, 15, 6, 20, 10, -17, -8, -4, -3, -18, -32, -49, -45, -43, -38, -43, -21, -44, 2, -16, -7, -6, -8, 1, 24, 4, 3, -14, -15, 4, 22, 0, -7, -11, 14, 3, -6, -5, -37, -7, -37, -10, -36, -40, -35, -24, -20, -28, 0, -29, -13, -23, 11, -14, -26, -37, -63, -4, 15, 7, 15, 10, -9, -8, 6, -9, -27, 6, 2, 6, -49, -42, -43, -46, -35, -39, -28, -47, -37, -24, -19, -59, -68, -60, -54, -34, 0, 8, 5, 18, 8, -18, 18, -16, 32, 43, 51, 11, -18, -3, -7, -29, -48, -71, -43, -45, -39, -77, -41, -47, -71, -72, -26, -41, -22, 1, 0, 17, 12, 12, 7, -2, 42, 87, 67, 66, 50, 41, 36, 4, 2, -22, -38, -43, -56, -70, -58, -71, -83, -66, -61, -51, 13, 6, -6, 12, -7, 5, -8, 11, 85, 44, 52, 109, 114, 76, 50, 37, 45, 34, 22, -10, -10, -45, -74, -79, -81, -61, -55, -40, -38, -17, 1, 2, -6, 12, 10, 14, 53, -11, 31, 50, 64, 88, 44, 78, 47, 79, 38, 26, -35, -5, -29, -1, -45, -44, -27, -19, -25, 0, 7, -5, 9, -7, 46, 11, 28, -8, -11, 15, 1, 42, 45, 56, 49, 64, 79, 19, 25, 47, 37, 11, -25, -7, -28, -23, 12, 5, 8, -15, 14, 13, 23, 15, 2, 26, 17, 6, -7, 11, -19, 28, 15, 55, 37, 38, 28, 36, 44, 1, -2, -3, -7, -14, 6, 11, 15, -18, 5, 2, -13, -23, 32, 53, 30, -31, -21, -18, -21, -11, 9, 32, 21, 11, 26, 32, 27, 14, -2, -20, -29, -15, 10, 20, -4, 15, -9, 1, -4, -5, -7, 11, 12, 0, -20, -4, 4, -26, -18, 25, 10, -1, 43, 23, 44, -1, 35, -4, -18, 0, 11, 47, 15, 19, 19, -2, 4, -57, 12, 38, -5, -2, 0, -6, -4, 4, -12, -5, 2, 33, 55, 48, 16, 34, 35, 14, -10, -31, -9, 59, -17, 19, 1, -1, -24, -66, -18, -49, -57, -25, -2, -39, -12, -29, -22, 1, -16, 16, 16, 0, 25, 24, 7, 15, -14, -35, 10, 28, 8, -5, -1, 17, -35, -20, -50, -31, -9, -19, 3, -33, -9, -20, -4, -4, 19, 20, 32, -4, -12, 16, 19, 40, 22, 0, 12, 40, 3, 18, 4, -2, -50, -38, -49, -44, -35, -27, -26, -16, 14, -19, -23, 10, 4, 6, -4, 12, 12, 37, 52, 13, 3, -42, 10, 18, -17, 19, -3, -13, -16, -10, -13, -35, -32, -67, -63, -9, -9, -23, -25, -26, -10, -3, 7, 9, 7, 19, 55, 19, 10, -8, -21, -4, -16, 4, -10, 1, -18, 21, 10, -3, -43, -37, -61, -74, -50, -48, -49, -31, -10, 10, -14, 7, 21, 20, 4, -3, 52, 14, -12, 1, 19, -14, 9, 7, 4, 14, 27, 13, -37, -32, -17, -37, -36, -24, -20, -44, -3, -15, -27, 3, 1, 27, 1, 17, 70, 14, -17, 10, 13, 18, -13, -3, -6, 14, 12, 8, -5, -18, -33, 16, 62, 51, 10, -40, -17, 16, -27, -12, 5, -25, -19, -14, -10, 24, -4, 4),
  9 => (-14, 10, -12, 16, 12, 7, 18, 13, -8, -8, -11, 10, 19, -12, -14, 11, 17, 15, 11, 11, -9, 15, 1, -10, 10, -7, -4, 13, 10, 2, -10, -11, -1, 7, 12, 12, 12, -6, -12, -14, -18, 12, 19, -16, 17, 5, -17, 2, -3, 14, -6, 5, -14, -10, 10, 12, 11, -8, 19, -20, 1, -15, 2, 1, -15, -9, -12, -17, -18, 0, -4, 5, -21, -30, -17, -5, -6, -23, -11, 9, 14, 0, 11, 19, 10, -10, 12, 6, -6, 4, -3, 12, 10, 2, 9, 0, -1, -20, -41, -19, 2, -11, -35, 20, 11, -3, 15, -16, 7, 12, 18, 10, -20, 2, 7, -3, -6, 12, -19, -8, 13, 3, -6, -5, -1, -17, -15, -33, -55, -32, -49, -47, 12, 10, 16, -1, 17, 2, 12, -14, 17, -5, -3, 9, -12, 3, 6, -8, -18, -16, -11, -36, -28, -33, -49, -29, -10, -9, 7, -30, -21, 19, -17, -6, -21, 14, -10, 12, 15, -16, -7, 0, -3, -5, -4, -13, -1, -31, -32, 22, 25, -39, -50, -55, -31, -22, 0, 11, 9, 0, -18, 9, -23, -14, -17, 10, -3, 15, 20, 7, -6, 11, -1, -22, -6, -48, -43, -11, 17, -43, -32, -34, -35, -44, -26, 18, 5, -20, -10, 2, -10, 4, 6, 20, 7, 17, 19, -12, 10, 7, 15, -5, -53, -17, 23, 7, 32, -29, -36, -47, -41, -24, -39, -27, -22, -2, -13, 21, 4, -4, -18, -15, -20, 1, 2, -21, -8, 16, 5, -41, 14, 26, 34, 63, -2, -29, -47, -45, -51, -25, -49, -30, -45, -1, -17, 15, -5, 9, 19, -2, -7, 10, 2, -11, 18, -10, -14, -8, 8, 39, 0, -1, -8, -5, -42, -23, -30, -38, -64, -12, -23, -19, 3, 16, 12, 0, -21, 1, -1, 12, 9, 13, 7, -9, -41, 12, 9, 12, 13, 7, -36, 4, -23, -15, -66, -22, -40, -58, -24, -40, 15, 14, -14, 2, -7, -7, 19, 12, -12, 18, 20, -7, -26, 6, -23, -18, -1, -23, -14, -43, -6, -7, -9, -11, -53, -35, -51, -23, 3, 7, -9, 10, -7, 3, 19, -1, 6, -19, 0, -18, -29, -87, -40, -42, -47, -25, -42, -30, -38, 19, -1, 14, -8, -23, -37, -35, -11, -10, -6, 16, -11, 7, 11, 1, 20, -21, 7, -15, -42, -83, -54, -43, -32, -29, -30, -37, -38, 8, -16, 15, -1, -28, -40, -21, 9, -16, -6, 10, -5, -9, -14, -12, -15, 18, 6, -6, -20, -32, -28, -10, -33, -7, -28, -44, -9, -22, -31, -7, 14, -9, -32, -24, -11, 14, -31, -18, -13, -12, -13, -20, -10, -2, -14, 6, -15, 1, 24, 14, -9, 20, -23, -44, -26, -10, -26, -25, -1, -48, -28, -21, -8, -14, -25, -3, -8, -8, -11, -5, 15, 14, 22, 11, 15, 30, 13, -1, 23, 50, 13, 0, -13, 9, -15, -13, 18, -6, -31, 6, -19, -11, -17, -7, -7, -2, 1, 20, -12, -15, 2, -12, -14, 27, 35, 20, 39, 57, 30, 58, 12, 14, 22, 0, -12, -4, 2, -27, -36, -2, -12, -10, -4, -8, 13, 20, 7, 6, 5, -12, 12, 14, 13, 17, 64, 25, 45, 23, 13, 34, 38, 30, 34, 7, 32, 29, 13, 21, 31, 6, -6, 0, 5, 3, 2, -8, 27, 28, 61, 43, 38, 7, 15, 1, -6, 14, 23, -10, 5, 11, 26, 11, 29, 29, 3, -5, 27, 1, -12, 1, -17, -1, 10, 6, 12, 32, 53, 56, -3, 31, -4, -28, -14, 15, 32, 13, 23, -3, 13, 27, 5, 30, 25, -37, -14, 13, -12, 0, 0, -3, -18, 9, 36, 3, -21, 8, 0, -15, -57, -27, -61, -14, -18, 24, -8, -8, 13, 7, -19, -26, 21, -4, -9, -27, -20, 1, 9, 18, -20, 8, 11, -7, -15, -6, -8, -51, -37, -36, -52, -35, -36, 3, -20, 15, 27, 10, -1, -56, -25, -10, 16, -3, -22, -1, -7, -15, -18, -21, -15, -17, 7, -5, -10, -56, -65, -39, -45, -24, -27, 3, -46, -15, 1, 21, -3, -9, -32, -24, -4, -29, -27, 19, 2, -16, -16, 20, 10, -36, -18, -14, -5, -48, -46, -64, -52, -32, -16, -17, -5, -21, -24, 8, -17, 0, -36, 1, -21, -5, 9, 15, -9, -6, -7, 6, -16, -9, -21, -22, -20, -27, -24, -41, -36, 1, -32, -15, 0, -9, -4, -3, -20, -38, -21, -30, 3, 17, -18, 22, -2, -13, -16, 13, -19, -12, 9, -42, 1, -16, 17, -3, 8, -20, -12, -30, -5, -2, -17, -9, -11, -26, -41, -19, 23, 15, 0, 3),
  10 => (20, 5, 8, -12, 4, -12, 19, -17, 18, 9, -6, 17, 13, -14, 4, -48, -24, -22, 8, -16, 11, -13, 7, 14, 11, -5, -18, 6, 7, 3, 12, 15, 16, 1, -19, -15, -3, 15, 7, -16, -13, -42, -8, -28, -34, -4, 17, -7, -50, -26, -27, 18, -14, -5, 17, 16, 15, 12, -5, 9, -13, -2, 4, 17, 21, 0, -11, -10, 23, 47, -5, -35, -66, -20, 62, 63, -19, -63, -65, 7, -12, 10, -20, 1, 2, 13, -16, 5, -1, 16, -12, 17, 16, 31, 8, 52, 6, -25, -44, -24, -21, 31, -5, -16, 16, -25, -63, -12, 26, 15, 7, 10, 19, 9, -7, -6, -13, 4, 0, -14, 33, -21, -13, -19, -54, -81, -8, 73, 27, 5, 6, 24, 30, -32, -42, -29, 12, -15, -9, -2, -18, 4, -14, 15, 1, 3, 7, 18, 21, 31, -8, -66, -103, -71, 14, 56, 62, 39, 10, 20, -7, -26, -15, -42, -22, -24, -16, 17, 15, -1, 0, -7, -10, 8, 13, 26, 85, 48, -37, -117, -128, -49, 25, 50, 38, 12, 23, -9, -22, -28, 13, -11, -39, -68, 3, 1, 14, 11, -17, -5, 19, -7, -8, 75, 60, 41, -76, -85, -118, 4, 46, 42, 51, 56, -26, -32, -15, -34, 17, -10, -58, -46, -12, -4, 9, -20, -14, -3, 7, -19, -38, 22, 69, 1, -66, -118, -95, 17, 71, 59, 46, 34, -31, -84, -43, -21, -19, -19, -25, -34, -57, -39, 14, 10, 20, -16, 2, -6, 1, 51, 16, -37, -88, -111, -28, 26, 59, 33, 28, 0, -40, -38, -55, -19, -1, 5, 14, -54, -29, -22, -16, -9, -20, 10, -17, 11, 0, 47, 11, -60, -103, -73, -30, 13, 52, 31, 32, -2, -1, -42, -44, -11, 18, 24, 17, -22, -31, 33, 9, 12, 18, 10, 2, 35, 39, 41, -8, -36, -116, -86, -16, -11, 70, 54, 18, -2, -33, -49, -19, -5, -6, 47, 24, -1, 1, -22, 16, 1, -4, 3, 10, 38, 18, -21, -7, -68, -90, -33, 28, 27, 37, 34, -28, -14, -42, -41, -23, -38, 0, 26, 19, 1, 10, -59, 10, -1, 6, -9, -2, 32, 52, -11, -70, -79, -80, -8, 34, 3, 40, -6, -27, -58, -28, -35, -7, -17, 10, -11, -8, 21, -35, -43, -14, -4, -3, -3, -3, -4, 63, 13, -72, -119, -52, 6, -22, -10, 14, -18, -28, -58, -33, 2, 20, 5, 44, -17, 4, -1, -19, -34, 11, -16, -18, 3, -11, 35, 41, -33, -79, -56, -35, -29, 3, -15, -1, -5, -12, 8, -26, -5, 12, 23, 41, 9, -5, -52, -60, -50, -18, 10, -5, -14, -53, 37, 37, -22, -63, -25, -5, 3, 8, -6, 0, -1, -25, -36, -40, 2, 5, -6, 24, 1, -34, -50, -65, -51, 9, -9, 19, -10, 7, 45, 44, -22, -30, -22, -28, 28, 36, 13, 1, 8, -41, -13, -12, -27, -1, 23, -3, -22, -37, -64, -48, -42, -11, 16, -3, -18, -29, 4, 43, 2, -34, -12, -12, 27, 22, 8, -25, 2, -25, -47, 2, 1, -1, -28, 34, 3, -91, -73, -54, -11, 20, -18, -15, 2, -29, 17, 11, 2, -25, 1, 3, -5, 12, 9, 21, 32, 1, -13, -9, -6, 2, 5, 14, -39, -41, -44, -72, 9, 19, -18, -9, -13, -14, 6, 44, 20, 7, 23, 18, 5, 15, 13, 11, 24, -9, 10, -9, 4, 12, 14, -11, -30, -58, -40, -42, -9, -12, -8, -11, 12, 13, 8, 11, 13, 3, 27, 21, 31, 23, -12, 25, 40, 38, 10, 17, 3, -21, -19, -4, -27, -23, 3, 30, 36, 10, 11, 18, -15, 5, -9, -12, -16, -10, 26, 33, 17, 1, 37, 16, 29, 12, -31, 20, 4, 27, -19, -6, -36, -30, -12, 22, 34, 4, -5, -18, 14, -2, 4, -15, -22, 5, -11, 5, 18, 7, 2, 21, -4, 20, -16, -23, 21, 27, 17, -9, -9, -7, -34, -20, -7, -17, -15, -13, 3, -25, -4, -4, -6, 2, -5, -1, 7, 2, 41, 16, 8, -9, -12, -8, -16, 8, -6, -11, 38, -5, -13, 0, 8, -3, 10, 13, 5, -4, -21, -2, -5, 17, 5, -25, -12, -33, 3, 13, -5, 30, 1, -13, -1, 4, -26, -16, -16, 43, 7, 5, -9, 2, 18, -13, -2, -11, 2, -27, -22, -25, 4, 3, -41, -18, -9, 0, 14, 23, 16, -5, -34, -23, -17, -37, -29, 6, -7, 12, -6, -3, 5, -8, 5, -15, -7, 14, -15, -18, -8, -49, -3, -34, 17, -27, -17, -10, 0, 13, 6, -8, -72, -37, -47, -27, -3, -10, -8),
  11 => (-18, 5, -4, -2, -2, 15, -5, -8, -18, 5, -14, -8, 10, -13, 10, 33, 61, 29, -36, -24, -2, 3, 18, -16, -5, 20, -14, 12, -15, 11, -12, -14, -6, -9, -17, -14, -6, -13, 14, -38, -46, -28, -21, 24, 49, 60, 33, -14, 19, 22, 66, 8, 10, 13, 17, 17, -4, 19, 8, -19, 18, -11, -19, -12, 15, -1, -21, -66, -22, 15, 36, 50, 34, 12, 0, -14, 0, 9, 67, 53, 5, 26, -12, -16, 8, -14, 5, 14, 9, 15, -20, -18, -5, -23, -28, -41, 34, 30, 33, 39, 10, -8, -15, -2, 0, 10, 16, 5, -40, -11, 15, -2, -19, -7, 11, 12, -6, -9, 15, 10, -29, -52, -43, 7, 20, 34, 4, 8, 35, -8, 20, 5, 4, 10, 14, 13, -28, 8, -3, 9, 20, 7, -16, -5, -10, 0, 2, 4, -77, -113, -10, 40, 18, -2, -4, 27, 8, -24, 10, -1, -6, 20, 47, 47, -42, 5, 12, -14, -16, 3, -3, -13, -15, -6, -15, -6, -101, -47, -20, 24, 41, -4, -23, 12, 18, -2, -15, 0, 8, 16, 37, 25, 13, -17, -7, -16, -17, 18, 9, 17, 6, -11, -28, -59, -93, -12, 30, 15, -13, 0, -62, -7, 13, -14, 13, -4, 5, 4, -38, 38, 23, 1, -7, -12, 12, -13, -5, 15, -19, -9, 1, -29, -45, 8, 37, 39, 23, -51, -43, 7, -8, -12, -33, -13, -20, -31, -17, 33, 30, 36, 4, -16, 2, 20, 17, 2, -15, -11, -3, 3, -40, 23, 38, 46, -13, -51, -37, -4, 3, -14, -9, -22, -40, -21, -2, -12, 29, 3, -34, 1, 18, -6, 7, -20, 10, 17, -26, -44, 16, 11, 54, 52, -43, -58, -57, 7, -14, -2, -3, -5, -18, -39, -36, -11, 4, 42, -17, -10, -14, -19, -4, -4, -7, -26, -33, -72, 35, 17, 66, 15, -79, -74, -50, 1, 0, 4, -15, -18, -18, -21, -46, -24, -17, 23, 0, 9, -10, 18, 3, -5, -14, -10, -3, -17, 59, 48, 55, 5, -78, -11, 3, 20, -2, -35, -13, -50, -32, -16, -26, -22, -7, 5, -2, 13, -15, -14, -14, 11, -1, -13, -43, 11, 83, 69, 49, -3, -78, 2, 5, 17, -3, -16, -48, -65, -69, 1, -15, 1, -35, 7, 0, 10, 9, -2, 4, 19, 40, -25, -64, 17, 55, 22, 12, -43, -95, -22, -9, 33, -1, -2, -43, -99, -70, -13, -9, -2, -40, -21, -25, -7, 8, 10, 14, -7, -19, -73, -63, 13, 43, 17, -12, -38, -53, -12, 38, 41, 16, 14, -31, -75, -62, 5, 30, -18, -39, -3, 19, -52, -19, -14, 1, 3, -5, -50, -48, 34, 3, 22, -7, -13, -55, 2, 22, 68, 39, 55, -40, -23, -15, -14, 7, 1, -24, 8, 29, -20, -6, 19, 5, -4, -15, -57, -41, 15, 15, -8, 15, -41, -58, 26, 38, 36, 51, 15, -56, -12, 27, 28, 24, 30, 11, 37, 35, -14, 8, 0, 14, -9, -6, -40, -40, 0, 29, -28, -22, -15, -53, 17, 44, 45, 51, 21, -50, -70, -35, -8, 19, 21, 8, 51, 76, -21, -12, 6, -9, 16, -10, -57, -42, 9, 13, -20, -34, -54, -42, 9, 40, 62, 43, 13, -28, -18, -50, 35, 40, 44, 12, 45, 35, -7, -6, -3, -15, -1, 5, -77, -4, 8, 3, -51, -50, -66, -35, -4, 45, -1, 23, 10, -9, -18, 4, 27, 29, 16, 31, 58, 30, -65, 5, -12, -6, -16, -6, -76, -31, -13, -27, -41, -51, -58, -18, -13, 13, 12, 4, 28, -38, -16, -6, 20, 25, 42, 26, 40, 42, -34, 16, -13, 2, -19, 21, -45, -51, 4, -42, -40, -73, -67, -21, 4, 26, 17, 38, 34, 4, 20, 2, 24, 34, 50, 32, 38, 21, -35, 12, -10, 9, -7, 15, -32, -47, -8, -46, -49, -56, -72, -57, -8, 39, 13, 36, 2, -12, -28, 19, 22, 30, 16, 42, 26, 20, -41, 4, 2, -19, -7, 0, -1, -30, -3, -31, -62, -49, -55, -10, -41, 36, -10, 18, 8, -18, -8, 4, 3, 18, 20, 36, 15, -14, -62, -13, -16, 16, 11, -13, -38, -48, -37, -43, -22, -31, -15, -13, -8, 4, 12, 19, 15, -35, -2, -22, -15, -14, 11, 23, 18, -46, -45, 0, 8, 18, -1, -5, -18, -54, -50, -9, -8, 10, 18, 10, 9, -7, 27, 25, 1, -10, 2, 6, 7, 11, 11, 7, -6, 3, -3, -9, 6, 8, 9, 11, -17, 1, -12, -2, -18, -5, -9, 21, 18, 26, 11, 47, -8, 2, -3, -22, -8, 7, 37, 35, 6, 7, -1),
  12 => (-10, 1, 8, 9, 14, 17, 18, 0, -8, 11, 8, 5, -13, 1, -11, -11, 17, 12, 7, 10, -24, -2, 6, 9, -3, -19, 16, 6, -19, -8, 6, 13, 17, -20, -17, -15, -11, -19, 4, -14, -1, -19, -27, -11, -15, -40, -57, -47, -36, -19, -23, 22, -3, -6, -9, -19, 18, 4, 7, 6, -18, -4, -4, 2, 6, 23, 20, -26, -4, -4, -24, -49, -34, -20, -56, -20, -16, -14, 2, 0, 15, 26, 8, -19, 8, 15, 5, -1, -13, -19, 3, -10, -15, 4, -37, -19, -3, 7, -9, -22, -7, -25, -35, -36, -5, -16, -8, 13, 3, 20, 9, -14, -2, 9, 3, 14, 18, 4, 1, 13, 11, 27, 6, 20, -12, 9, -24, -43, -27, -22, 6, 17, -23, -31, -58, -16, 2, -21, 9, 13, -10, 7, -2, 9, 7, -5, -13, -14, 42, 18, -1, -32, -32, -26, -18, -7, -3, 0, -7, -25, -5, -1, -31, -17, 22, -10, -17, -19, -16, 2, 17, 6, 2, -11, -3, -46, 17, 43, 67, 25, 45, -8, -3, -25, 21, 18, 31, 18, 3, 9, 5, 27, 12, 19, 20, 8, 0, 13, -14, 17, -14, -11, -31, 5, 24, 57, 35, 27, 33, 36, 3, 24, 11, 29, 56, 38, 41, 9, 35, 27, 25, -26, -18, 1, 10, -10, -11, -11, 1, -7, 9, 34, 44, 48, 17, -11, 11, 30, 19, 31, 25, -6, 37, 57, 38, 51, 22, 45, 13, 4, -5, 16, 13, 7, 16, -15, 8, -13, 4, 51, 46, -55, -23, -39, -9, 8, 26, 16, 19, 23, 17, 26, 58, 59, 54, 42, 45, 57, 18, -2, -16, 9, 8, -18, -16, -2, -17, -3, -27, -78, -76, -72, -101, -57, -35, -91, -43, -23, -7, -31, -28, 0, -4, -18, -3, 54, -11, -14, -5, -1, -11, -10, 2, 16, -16, -20, -25, -56, -77, -73, -75, -43, -70, -78, -58, -76, -83, -101, -48, -59, -52, -68, -38, 36, 8, 5, 20, -19, 2, -17, 13, -19, -43, -25, -9, -20, 9, -4, -20, -49, -53, -61, -56, -67, -76, -81, -61, -63, -76, -72, -66, -25, 30, -8, -12, -5, 4, 16, -7, 0, 4, 42, 44, 31, 56, 67, 17, 15, 38, 30, 29, -9, -3, 19, -27, -7, -31, -40, -55, -38, 0, -38, 3, -3, 5, 10, -3, 6, -12, -3, 1, -2, 23, 38, 51, 38, 42, 28, 33, 25, 4, -14, 17, 31, -5, 13, -71, -91, -66, -35, -14, 1, 5, -9, 6, -16, 27, -1, -19, -7, -10, -7, 12, -9, 33, 34, 19, 14, 37, 34, 34, 27, 21, 15, 3, -25, -48, -8, -1, -20, -17, 10, 31, 1, 7, -66, -64, -12, 7, 21, -12, -11, -12, 26, 23, 36, 25, 16, 59, 16, 22, 8, 21, -6, -19, 11, 5, 8, -8, 3, 29, 0, -17, -38, -39, -7, -14, 4, 11, -43, -2, -16, -19, -28, 20, 4, 18, 35, -16, -32, 11, -12, -28, 6, 14, 18, 17, -2, -43, -45, -35, -18, -41, -41, -19, 48, 33, -19, -6, -5, -8, -1, -9, 9, -1, 23, -13, -43, 32, 24, 4, -17, -6, 19, -17, 7, -53, -42, -23, -5, 12, 33, 52, 8, 30, 9, 3, 6, -6, 17, 22, 10, 18, 15, -14, -27, 15, 54, 36, 19, 1, 2, 16, -1, 18, 6, -39, -6, -5, 26, 73, 42, 4, 21, 20, 11, -6, 20, 22, -9, -20, 2, -5, -18, -8, 16, 25, -3, -19, 13, -8, 18, 39, 6, -15, -26, -21, -8, 16, 10, 23, -3, 8, -12, -4, -1, 2, -14, -15, -48, -30, -40, -13, 11, 20, -1, 20, 1, 12, 3, 25, -31, -23, -3, -16, 1, -18, 10, -14, -3, -6, -13, -19, -10, 14, -23, -3, 22, 2, 6, -8, -4, -4, 0, 20, -8, 14, 2, -14, -17, 8, -7, 2, 5, 13, 9, -5, 5, 13, -24, 5, -20, -11, 35, 8, 20, -19, -15, -7, -17, 1, -7, 2, -19, 4, -20, 6, -18, 23, -3, -27, -2, -19, -31, -30, -22, -48, -35, -16, -8, -10, -20, 8, -14, -7, -18, -1, -37, -6, -6, -4, -4, 4, -3, 9, 3, 4, 10, 8, -6, 3, -20, -5, -30, -10, -12, -25, -37, -43, -2, 6, 3, 32, 21, 16, -7, -11, -6, -18, 0, -9, -19, 14, 4, 17, 25, -4, 2, -33, -21, -1, -4, -14, 14, -20, -22, -18, -66, -31, -25, 9, 11, 45, 26, 35, 5, 9, 8, -16, -12, 18, 19, 13, 4, -8, 22, -14, 24, 33, 51, 21, -39, -8, 48, 42, 8, -13, -30, 32, 42, 25, 36, 42, 1),
  13 => (19, -4, 9, 15, -13, -17, 4, 10, -16, -1, 12, 0, 3, 14, 20, -1, -20, -8, 24, -13, -14, 10, 20, 2, 13, 8, -1, 9, 6, 2, -13, -4, 3, -1, 14, 6, 16, 5, 52, 59, 33, 38, 23, 12, 15, -9, 21, 38, -9, -17, 7, -3, -6, -12, 3, 15, -19, -6, -6, -16, -15, -12, -14, 2, -9, 82, 36, 9, -8, -17, -15, 10, -15, 20, 40, 25, -8, -15, -2, -9, -18, 10, -14, 2, -3, -18, 7, -4, -2, 13, -16, 10, 52, 23, -37, 3, -11, 33, 54, 10, -21, -9, 3, -26, 0, -20, 13, -13, -16, 13, 2, 16, -7, 12, 9, -15, 0, -7, 6, 7, -14, -57, -9, -32, 21, 50, 31, -9, -58, -23, -33, -35, -21, -11, 18, -17, 0, -15, 9, 18, 11, -3, 5, 14, -15, 1, 1, -17, -20, -27, 14, 35, 36, 14, -47, -61, -59, -44, -35, -46, -11, 18, 23, -6, -12, -2, 1, 6, -5, 15, -16, 15, -13, 0, 15, -2, 7, -4, -8, 40, 44, 6, -57, -47, -58, -76, -6, -32, -22, -3, -8, -14, -13, -14, 3, 11, 2, -16, 3, 14, 0, -2, -2, 3, 0, 22, 43, 28, 11, 4, -27, -10, -17, -26, -37, -45, -2, 11, -1, 0, -1, 6, -17, -7, -18, -19, -10, -14, -7, 12, 34, 2, 19, -13, 4, 1, 12, -17, -40, -18, -30, -58, -50, -26, 9, -11, 3, -12, -4, -20, 7, 19, -11, -18, 0, 16, -2, 18, 26, -4, 11, -21, -26, -3, -4, -6, -24, 9, -33, -31, -30, 41, -21, 6, 11, -6, 10, 0, 14, -6, 19, 4, -2, -11, -13, -16, 15, 55, 9, -7, -5, 17, 7, 22, -21, -10, -13, 16, 5, -1, 44, 28, -19, -36, -5, -9, 19, 13, 12, -7, 19, -13, 11, -44, -7, 13, 28, -6, -22, -16, 12, -7, -10, -25, 9, -10, 26, -2, 24, 39, 17, -34, -17, 8, -9, -9, -3, 14, 4, 6, 1, -24, -23, -11, 19, -4, 6, -50, -20, -71, -38, -43, -29, -1, 3, 35, 16, 6, 6, -26, -1, -24, -2, -3, 12, -6, 6, 9, -6, -75, -34, -12, 22, 50, 12, -39, -38, -46, -48, -124, -68, -60, -37, -47, -18, -4, -27, -23, 11, -20, 1, -20, -3, 4, -4, 17, -30, -83, -58, 12, 38, 44, 31, 30, 13, -22, -54, -104, -115, -114, -100, -109, -113, -72, -64, -54, 9, -3, 3, 1, 20, 13, -15, -9, -28, -55, -27, 21, 24, 10, 29, 35, 10, 20, -12, -32, -61, -77, -96, -102, -90, -70, -57, -77, -20, 2, 10, 8, 11, 0, -18, 15, -25, -39, -40, 13, 29, 12, 0, 16, 35, -5, 6, 8, -19, -21, -60, -82, -68, -54, -46, -54, -52, -25, -8, 9, 18, -19, 19, -8, -15, -66, 17, 22, 10, -23, 1, 9, 1, -2, 11, -15, -10, 0, -7, -32, -27, -19, -26, -59, -48, -11, 25, 4, 17, -19, -10, 8, -4, -111, -20, 17, -3, 5, -8, 32, 6, -18, 9, -12, -1, 16, -27, -26, -6, 5, 12, -20, -71, -4, -18, 4, -11, 16, -20, -10, -50, -92, -38, 4, -2, 29, 24, 29, 8, -13, 20, -8, -8, 39, 24, -2, 30, 31, 2, 17, -23, -8, 12, 5, 16, -17, 6, -7, -19, -65, 5, -21, 41, 31, 17, 9, 8, -11, -6, -22, 7, 24, -6, 19, 16, 12, 14, 24, 19, 11, -6, -2, -20, -15, -19, 13, -22, -26, 6, 9, 13, 36, 43, 32, 16, 8, 16, 2, 7, -4, 29, 15, 13, 35, 25, 4, 18, -20, 3, 5, 18, 5, -5, 1, -19, -31, -25, -20, 24, 2, 17, 30, 5, 26, 6, 36, 51, 27, 31, 55, 14, 17, 25, 38, 19, 12, -6, -13, -2, 8, -2, -11, -44, -59, 0, 14, 18, 39, 40, 13, 5, -6, 13, -4, 6, 5, 49, 66, 24, 25, 21, 17, 29, 19, 4, -20, 8, 2, -10, -9, -65, -36, 13, -22, 9, 32, 33, 23, -9, -2, 28, 18, 17, 55, 59, 61, 14, 13, 2, 37, 3, 13, 45, -60, -5, -7, 15, -17, -48, -25, -7, -27, 20, 37, 55, 41, 21, 24, -1, 23, 28, 19, 29, 46, 73, 46, 39, 44, 17, 22, -18, -20, 19, -12, -15, -14, -51, -26, -8, 14, -12, 37, 39, -4, -20, -1, 13, 2, 9, 6, 27, 48, 5, 14, 10, 31, 39, -11, -21, -6, 5, -2, -7, 20, -13, 18, -12, 36, -5, 12, 15, 11, -1, -16, -13, 16, 7, 25, 14, -1, -4, -15, 25, 23, 20, -13, -33, 13),
  14 => (5, -17, -16, -13, 20, 18, -16, -17, 14, 3, 1, -7, 4, 17, 18, -31, -18, -11, -56, -49, -13, 20, -3, -8, -4, 7, -19, 6, 11, -3, -19, -5, -13, -4, 18, 10, 4, 14, 47, 39, 29, 10, 55, 6, 40, 26, 25, 45, 17, 23, 40, 21, -12, 13, -20, 12, 5, -6, 19, -15, 1, -4, 18, 1, 11, 54, 28, 71, 43, 59, 64, 42, 60, 48, 73, 66, 51, 30, 13, 17, 7, 13, 7, 8, -6, 16, 10, -7, 14, 8, 20, 11, 39, 47, 54, 35, 21, 40, 82, 14, 31, 0, -9, -27, 11, 1, 4, 4, -28, 4, -12, -9, 6, 18, 7, -16, -1, -19, 11, -3, 2, -38, -30, -20, -30, 34, 58, 23, 22, -1, 4, -6, -12, -12, -27, -24, -8, -1, -17, 5, -8, -14, -15, 9, 6, -4, -6, 40, -4, -73, -94, -25, 8, 44, 36, 17, -3, -9, 8, 41, 13, -15, -36, -27, -28, -10, 19, 19, 12, -8, -8, 20, -11, 3, -20, 39, -13, -29, -16, -4, 61, 47, 43, 34, 22, 14, 47, 22, 53, 17, -14, -36, -15, -58, -13, 20, 11, 6, 2, -15, -16, 8, -11, 63, -9, 10, 33, 3, 25, 32, 16, 21, 11, 24, 25, 25, 20, 0, -8, -57, -3, -39, -35, -21, 4, -7, -4, -18, 10, 0, 21, 35, 5, 9, 4, 9, 28, 32, 38, 27, 29, 2, 3, -25, -47, -21, -73, -94, -48, -33, -43, -7, 19, -9, 20, 17, -11, -18, 30, -10, -3, -5, -18, 6, 18, 45, 59, 35, 30, 49, 33, -27, -27, -38, -82, -94, -25, -20, -39, -17, 7, 14, -3, 19, 12, -29, -26, -25, -6, -6, -8, 19, 19, 10, 27, 24, 4, 0, 9, -36, -24, -61, -51, -62, -31, -1, 1, 12, 10, -18, -12, -2, -8, -63, -66, -2, 4, 43, 56, 47, 29, 16, 13, 17, -7, -9, -37, 0, -40, -52, -34, -68, -41, 15, 35, -40, 7, -13, -7, 6, 23, -79, -24, 26, 20, 81, 43, 32, 62, 9, 24, 39, 9, -14, 24, 7, 9, -24, -60, -52, -44, 3, 31, -32, -5, -19, -15, -10, -14, -62, 27, 67, 58, 62, 68, 68, 52, 71, 27, 44, 48, 33, 20, 62, 28, 31, 24, 8, -17, 59, 31, -17, -12, -12, 15, -19, -19, -55, 11, 39, 40, 30, 54, 39, 24, 53, 40, 72, 52, 60, 42, 66, 65, 79, 68, 9, 55, 61, 44, 21, 9, 14, -19, 10, -22, -26, 22, 24, -16, 10, 23, 42, 65, 21, -9, 4, 26, 4, 35, 37, 35, 70, 36, 42, 28, 60, 52, -28, 2, 12, 14, -19, -36, -46, 10, 44, 2, 10, 30, 20, 15, -5, -36, 10, 5, 42, 8, -10, 35, 48, 28, 70, 60, 59, 47, -20, 12, -20, -13, -10, -11, -8, 29, 24, 28, 36, 17, 18, 14, -16, 18, 1, 10, 4, 12, 7, 51, 24, 51, 84, 73, 47, 60, 7, 5, 1, -18, -10, -11, -11, 16, 23, 2, 3, 28, 21, -3, 7, 6, 15, 10, 23, 29, 44, 51, 45, 85, 108, 51, 47, 63, -4, -18, 17, 8, -15, -9, 11, -9, -24, -2, 3, 15, 13, -3, -16, 2, 8, 3, 54, 10, 39, 74, 69, 51, 47, 15, 17, 42, -13, 0, 17, 19, -8, 31, 27, 28, -21, 18, 23, 16, 27, 10, 27, 48, 31, 55, 53, 29, 29, 54, 46, 15, 32, 15, 8, 21, -40, -13, -6, 4, -8, -15, -12, 15, 30, 12, 28, 67, 64, 22, 13, 41, 41, 49, 28, 27, 22, 40, 63, 36, 45, -20, -12, -20, -24, 20, 12, -11, 13, -39, 13, 23, 26, 17, -45, 10, 26, 23, 2, 32, 27, 54, 44, 26, 35, 40, 34, 26, 14, 10, -3, -24, -33, 13, -3, -11, -11, -31, -12, 17, 26, 2, -35, 25, 35, 15, -2, -2, 2, 32, 30, 16, 66, 53, 21, -7, -13, -5, -34, -7, -4, -7, -3, 7, 20, -13, -37, -8, -2, -20, -45, 9, 10, -4, 24, 3, 9, 18, 13, 19, 6, 22, 18, -42, -59, -4, -16, -11, 1, -9, -12, 17, 7, -40, -36, 16, 29, 3, -34, -13, 19, 4, 7, -6, 1, 20, 40, -9, 17, 1, 5, -16, -30, -19, 12, -8, -30, 16, -3, 17, 4, 6, 10, 17, -35, 34, 14, 29, 5, 13, -17, -29, -19, 8, 22, 10, -19, -6, 7, -9, -34, 8, 2, -35, -41, -5, 3, 20, -7, 13, 30, -8, 56, 73, 65, 34, 39, -1, 21, 47, 33, 29, 59, 39, 2, 13, 22, 20, 20, 23, -3, 12, -4),
  15 => (-5, -9, 18, -3, -10, -14, -20, -16, 16, 19, -20, 3, -15, 16, -45, -41, 22, -30, -8, -22, -21, -27, -7, 8, -20, 7, 5, -19, -13, 12, -21, -9, -4, -18, -1, 13, -14, -9, 26, 14, 18, 25, -1, 22, 5, 16, -6, -3, -5, 3, 20, 13, 21, 20, -8, 16, -9, -3, -3, 4, -2, 12, -19, 15, 3, 3, 13, 31, 7, 28, 16, 23, 14, 31, 22, 34, -17, -22, -36, 20, 23, 10, -13, -4, 20, 20, -13, 4, 4, 5, 4, 9, 0, -1, -5, -29, -17, 0, 33, 24, 21, 21, 2, 21, 20, -31, -10, -49, -8, -2, -12, 6, -1, 4, -9, 13, 2, 14, -15, -32, 30, -23, -11, -34, 23, 29, 48, 16, 1, -2, -8, -8, -26, -12, -11, -26, -24, -7, 9, -6, -5, 4, -2, 2, -13, 0, -9, 7, -1, 1, -35, -5, -7, 11, 24, 28, -19, 7, -8, -26, -16, -33, -24, -21, -13, 10, 1, 17, 0, 6, -1, -17, -4, 17, -23, 27, -1, 0, 30, 14, -11, -10, 10, 18, 19, -14, -16, -9, 21, 16, -16, -46, -17, 47, -2, 6, -20, -3, 14, 4, -7, 0, 4, 31, 35, 35, 45, 20, -23, -3, -8, 4, -19, -17, -47, 1, 3, 16, -38, -27, -7, 29, -4, 8, 7, -18, -16, 17, -4, -1, 38, 45, 40, 43, 43, 7, 18, -18, 5, -6, -20, -37, 6, -24, -15, -15, -17, -41, 23, 62, 7, 14, 13, 18, -9, 19, -20, 10, 31, 14, -4, 13, -7, -37, -5, 5, -23, -53, -54, -61, -9, -30, -15, -17, -30, -3, -1, 50, 30, 4, -13, -3, 9, 16, 5, 4, 32, -22, -32, -24, -29, -64, -34, 8, -43, -27, -1, -86, -51, -20, -26, -10, 5, 35, -10, 38, 13, -5, 5, -19, 6, 16, 1, -6, -12, -92, -66, -54, -19, -68, -10, -15, -29, -48, -38, -40, -47, -17, -40, 0, 26, 19, 19, 17, 15, -9, 17, 10, 3, -3, 8, 12, -36, -75, -54, -43, -57, -52, -17, -23, -63, -40, -41, -59, -16, -28, -35, 6, 6, 18, 24, 22, 42, 29, -15, 20, 15, -8, -17, 42, -14, -4, -3, -10, 23, 0, 14, 19, -4, 11, 18, -21, -16, 17, -12, 6, 26, 42, 19, 21, 73, 4, -16, -15, -7, 10, 53, 47, 53, 44, 75, 68, 29, 61, 49, 41, 71, 62, 50, 34, 21, 13, 10, 13, 5, 18, 0, -1, 39, 31, 20, -14, -15, 12, 26, 38, 61, 60, 86, 87, 56, 38, 51, 23, 55, 48, 35, 19, 14, 38, 22, 11, 18, 28, -17, 8, 12, 35, -17, 3, 11, 0, -1, 19, 14, 39, 16, 8, 22, 23, 54, 18, 51, 23, 46, 49, 17, 41, 14, 41, 14, 9, 21, -22, -3, 19, 16, 6, -17, 16, 39, 14, -19, -7, 7, 2, 3, 15, 31, 32, 11, 16, 47, 55, 40, 28, 38, 5, 4, 39, 44, 26, -16, 14, -1, 6, 8, -3, 21, -27, -46, 1, 42, 21, -9, 18, 28, 72, 24, 15, 46, 51, 45, 13, 58, 18, 8, 48, 18, 0, 37, 51, 9, 3, 15, 15, 7, 5, -22, -21, 5, -17, -36, -25, 10, 2, 27, -12, 16, 55, 27, 38, 36, 56, 21, 24, 25, 25, -2, 12, -20, 16, -19, 16, -12, -27, -12, -33, -46, -30, -55, -32, -41, -75, -60, -58, -46, -31, 10, 10, 27, 18, -2, 27, 21, 16, -14, 30, -20, -6, 19, 18, -14, -9, 9, -11, -33, -71, -107, -62, -63, -29, -82, -72, -62, -63, -35, -24, 2, -22, -22, -49, -27, -34, -19, 17, 0, 20, 5, 4, -2, -7, -18, -55, -60, -45, -72, -62, -54, -46, -52, -91, -63, -65, -33, -16, -38, -25, -42, -75, -108, -59, -38, 11, -5, 17, 7, 4, 18, -11, -29, -49, -25, -36, -45, -79, -52, -49, -79, -95, -89, -42, -28, -47, -33, -51, -40, -80, -69, -59, -20, 14, 6, -3, 20, 4, -1, -4, -12, -21, -16, -45, -7, -44, -23, -60, -73, -87, -97, -58, -24, -30, -64, -18, -13, -88, -104, -33, -14, 19, -3, 14, -17, -1, -1, 5, -19, -29, 2, -29, -21, -1, -31, -37, -62, -81, -67, -60, -28, -50, -62, -71, -24, -34, -78, -63, -3, 31, 19, -8, -17, -1, -10, 1, 11, 3, 2, -27, -5, -17, -52, -32, -37, -23, -41, -47, -27, -66, -24, -15, -47, -19, -21, -13, -17, -17, -8, 6, 14, 9, 9, 4, -2, 9, 3, 3, -23, -8, -13, -2, 3, -1, -21, 0, 1, 6, -45, -50, -25, -33, -22, -23, -5, 3),
  16 => (2, 0, 2, 2, 19, 8, -17, 15, 0, -15, -20, -15, -7, -11, -6, -31, -40, 18, -3, -39, -22, -11, -14, 3, 20, 3, 0, 1, -1, 10, 12, -9, 3, -1, -13, -1, -18, -16, -3, 5, 28, 28, 0, -5, -38, -16, -12, -24, -9, 2, -15, -13, 3, -18, -8, 13, -10, -3, -13, 5, -5, -4, 21, 11, 19, -2, 21, 40, 65, 63, 33, -2, -3, -53, -62, -43, -11, 11, 6, 4, 11, 9, -9, 7, 9, 20, 5, 8, 21, 2, -18, -6, 19, 2, 8, -13, 18, -22, -23, -14, -31, -42, -37, -46, 6, -39, -24, -17, -5, 19, 17, 9, -6, -16, -7, -15, 9, 8, -3, -16, 40, 35, -12, 12, 32, 25, 19, -13, -53, -65, -20, -25, -18, -35, -40, -61, -68, -7, -6, -20, -1, 7, 3, 18, 12, -1, -3, 14, 20, 25, 11, 10, 31, -15, -31, -42, -27, -30, 0, -15, -47, 5, 30, -24, -23, -50, -13, -15, -19, 5, 14, -16, -17, -19, -10, -21, 20, 16, 11, 9, -35, -82, -72, -58, -24, 14, 32, 37, 31, 56, 30, -7, -13, -20, 25, -15, -21, -17, -13, 16, 20, -3, 10, 17, 27, 30, -23, -27, -64, -63, -28, -35, 30, 55, 43, 48, 48, 50, -25, -17, -44, -4, 9, 6, -19, 3, -3, 11, 8, -17, -27, -13, -28, -37, -31, -64, -49, -2, 10, 9, 28, 46, 41, 19, 12, -10, -15, -67, -64, 3, -13, 23, -18, -12, 10, 6, -1, -19, -52, -50, -50, -65, -57, -38, 1, -29, -3, 11, 3, 35, 32, 0, 3, -21, -34, -49, -53, 1, 11, -7, 3, 12, 12, 0, -15, 19, -28, -115, -60, -37, -13, -14, 1, -11, 11, 8, 30, 12, 17, -27, -28, -32, -34, -66, -82, 9, -20, 30, -18, -16, 11, 20, 5, -32, -42, -61, 2, 9, -2, 14, -28, 29, 10, 10, 47, 36, 19, -22, -46, -61, -56, -22, -28, 35, 6, -7, 16, -10, 20, 1, 37, 6, -12, 4, 57, 68, 49, 38, 29, 41, 24, 12, -29, -50, -56, -50, -56, -28, -54, -46, -53, 0, -3, -12, -3, -20, 19, 12, 40, 4, 21, 70, 54, 47, 24, 18, 23, 23, -7, -24, -40, -44, -67, -46, -60, -36, -46, -30, 0, -13, 26, -35, -14, -10, 17, -12, 29, 48, 45, 35, 30, 44, 6, -17, -7, -9, -15, -16, -54, -21, -33, -61, -84, -50, -23, -16, 17, 33, 7, -2, 9, 19, 2, -11, 13, 65, 49, 33, 34, 30, 2, -10, -7, -22, -24, -6, 8, -55, -38, -58, -49, -61, -3, 42, 58, 47, 3, -7, -18, 11, -1, -19, 25, 53, 27, -19, 2, -4, -13, -27, -32, -44, -34, -31, -37, -30, -31, -6, -26, -25, 25, 41, 78, 68, 7, -9, -14, -2, -14, -9, -3, -15, -9, -56, 4, 13, -30, -1, -37, -53, -49, -47, -58, -60, -24, 29, 29, 36, 61, 49, 51, 33, 58, -8, 14, -3, 11, -3, -29, -32, -32, -53, -50, -11, -46, -45, -46, -66, -44, -47, -15, -5, 21, 51, 30, 26, 58, 76, 27, 60, 74, -45, 7, 7, 19, -15, -37, -33, -61, -51, -40, -49, -58, -62, -27, -20, -25, -23, 5, 31, 31, 49, 43, 12, 40, 68, 62, 63, 67, -24, 1, 3, -5, -17, -41, 4, -65, -23, -14, -17, -31, -14, -8, 18, 19, -3, 23, 24, 50, 22, 17, 10, 24, 23, 48, 25, 58, -26, -6, 12, -9, -17, -14, 33, -29, -10, 0, 11, 2, 53, 18, 52, 12, 1, 32, 9, 24, 16, 19, 2, -9, 31, 28, 7, 19, -9, -18, -7, -2, 20, 10, 28, -15, 20, 34, 19, 41, 35, 41, 80, 46, 12, 36, 6, 27, 27, 26, -21, 2, 15, -4, 11, 25, -33, 7, -19, 4, 2, 49, 53, -10, 1, 38, 28, 26, 21, 38, 47, 45, 14, 15, 21, 6, -12, 8, 7, -8, 21, 29, -10, -4, -46, 8, 9, 20, -9, 42, 35, 0, 1, 26, 3, 29, 11, 22, 17, 41, 10, 46, 38, 17, -21, 22, -7, 25, 23, -4, -61, -30, -13, -7, -20, -20, -14, 46, 2, 1, -2, 19, 25, 5, 40, 27, 28, 14, 8, 5, -25, -1, 11, -9, -17, -31, -11, -41, -46, 4, 38, -14, 17, 7, -2, 26, -19, -31, -22, 15, 17, -21, 5, 10, 5, -15, -12, 23, -1, -23, -4, -13, -47, -87, -78, -35, -23, 14, 56, -4, 5, 16, -6, 11, -21, -55, -18, -55, 25, 1, -6, -6, -7, -36, -8, 10, -19, -21, -37, -58, -65, -76, -30, -72, -23, 47, 39),
  17 => (4, -10, -8, 8, 1, 5, -15, -15, -5, 6, -17, 20, 3, 19, -18, 10, 51, 18, -14, 10, -40, -50, -17, -6, 21, 13, -13, -2, 5, -10, 18, 1, -19, -6, -20, 9, -13, 3, 25, -3, 13, 21, 38, 3, 43, 51, 32, -4, 33, 2, 3, 4, 11, 19, -15, 18, -19, -16, -12, 16, 6, 6, -2, 6, 1, -19, -20, -6, 29, 11, 21, -3, -3, -23, -14, -19, 9, -32, 3, 27, 29, -11, 2, -13, 0, -9, -2, 20, -12, 4, -17, -7, -27, -66, -49, -22, -19, -14, -41, -29, -3, -34, -10, 25, 22, -9, 8, 2, -8, 23, -3, -2, -18, 11, 4, -4, 11, 9, -2, -6, -62, -24, -32, 6, 12, 13, -15, 11, -7, 14, 6, 8, 13, 23, 2, -29, -17, -73, -5, 7, -15, -10, -19, 8, -5, -10, -23, -20, -2, -9, -7, 19, 25, 45, 32, 39, 40, 26, 26, 23, 38, 18, -24, -40, -70, -19, 1, -4, -7, 9, 15, 0, 0, 20, -27, -42, -14, 36, 15, 27, 43, 66, 20, -12, 42, 36, 31, 12, 57, 4, -25, -30, -9, 35, 27, 17, -11, 9, -10, -21, -11, -6, -45, -36, 21, 6, 24, 12, 37, 20, 17, 0, -2, 29, 5, 27, 12, 21, -33, -41, -44, 1, -27, -8, -20, 13, -1, 16, 19, -15, -17, 12, 52, 23, 17, -18, 15, 15, 3, -7, 25, 32, 35, 1, -12, 29, -21, 13, 21, 14, 15, -41, -15, 7, 4, -8, -1, -17, 1, 31, 28, 0, -24, 28, 58, 36, 6, 15, 5, 27, -16, -19, -2, -21, -17, 15, 15, 14, 9, 13, 21, 10, -3, -2, 3, 23, 39, 39, 32, -23, 6, 15, 31, 31, 13, 7, 30, 9, 1, -17, -37, -13, 11, 22, 34, -24, 4, 42, -16, 11, -20, 6, 9, 73, 35, 37, 29, 24, 54, 31, 24, 28, 6, 7, 15, 8, 18, -17, 5, -14, -31, -7, 25, 13, -36, 22, 5, -8, 4, -9, 2, 46, 8, 17, 12, 3, 11, 31, 59, 45, 17, 14, 29, 22, 27, 2, -5, -6, -44, -24, 30, -6, -45, 36, 13, 18, 1, -16, -54, 15, -19, -23, 0, 38, 35, 61, 40, 39, 37, 34, 9, 33, 31, -1, -28, -5, 30, 8, 42, 15, -20, 46, 3, -1, -5, -7, -22, -38, 2, -11, -18, -24, -34, -36, -61, -37, -17, -30, -25, -18, -17, 24, -7, 0, 38, 45, 29, 25, 32, 44, 13, -10, -9, 11, 16, 33, 5, -15, -34, -74, -107, -113, -120, -92, -52, -71, -83, -38, -36, 0, -10, 34, -10, 0, 24, 30, 44, 71, -10, -1, 11, 1, 25, 23, -49, -99, -102, -107, -82, -69, -87, -33, -19, -75, -39, -67, -59, -39, -65, -39, 3, -1, 24, -4, 29, 21, 19, -18, 13, 17, 0, -69, -95, -95, -91, -107, -99, -76, -35, -20, 12, -62, -39, -72, -23, -29, -60, -67, -20, 8, 16, 16, -19, 27, 15, 14, 14, -19, -23, -59, -78, -67, -66, -70, -63, -103, -56, -35, -19, -67, -44, -43, -32, -16, -69, -44, -42, -5, -3, 21, -10, 52, -1, -19, -12, -20, -1, -79, -66, -42, -61, -59, -55, -25, -8, 26, -20, -19, -14, -39, -39, -26, -17, -25, -30, -29, -4, 6, 38, 65, -7, -10, 20, 8, -41, -50, -48, -33, -3, 34, 13, 27, 30, 3, -5, 24, -6, -6, 18, -26, -24, -33, -38, -22, -9, 36, 52, 59, 2, 6, 3, -14, -21, -16, -13, 7, 8, 8, 43, 65, 59, 12, -6, 38, 20, 20, 19, -10, 11, -12, -25, -57, -45, 23, 67, 59, 8, 9, -4, -9, 26, 65, 10, 3, 13, 13, 12, 30, 42, 37, -9, 17, 25, 2, 34, 17, 25, 32, 2, 19, 8, -4, 4, 38, -15, -15, -1, 16, 42, 30, 11, 18, 12, 28, 28, 44, 39, -1, 19, 0, 15, 22, 10, 27, -7, -20, 20, 50, 40, 37, 9, 17, 2, 17, -20, 15, 36, 67, 17, 42, 4, 25, 16, 25, 14, -14, 11, 30, 19, 0, -10, -11, 27, 50, 65, 3, 35, 62, 26, 21, 1, -3, -11, -12, 66, 56, 68, 5, 25, 28, 34, 8, -4, -8, -1, -9, -40, -30, 10, 3, 28, 31, 44, 70, 53, 45, 35, 61, 18, -20, 11, -12, 39, 37, 36, 46, -6, -1, -7, 10, -7, 16, 5, 6, 4, 0, 4, -29, 2, -3, 30, 62, 82, 37, 16, 98, -4, -17, -5, -17, 17, 25, 30, 0, -9, 9, 29, 0, -9, -6, -8, 50, 23, 22, -4, -17, -19, 11, 36, 78, 54, 53, 42, 36),
  18 => (17, 13, -18, -15, -20, -5, -14, 8, 18, 13, -17, -14, 2, 13, 13, 11, -14, 2, -7, -12, -20, -18, -15, 8, 17, 20, -8, -4, -7, -15, 7, 19, 16, 7, 10, 7, -1, 11, 1, -2, 14, -13, -49, -11, -6, 10, 4, 10, -6, -9, -10, -17, -30, 3, -19, -9, -17, -16, 11, 7, -18, -16, 3, 20, 7, -19, -23, -6, -2, -6, 10, -4, 26, -29, -8, 11, 36, 20, 11, 11, 13, 0, 11, 17, 2, -16, 10, 11, 21, -18, -19, -6, -4, -14, -1, -39, 11, 1, -17, -35, -2, -6, -13, 0, 16, 9, -5, 44, 48, 25, 11, 0, -11, -1, -3, -7, 17, 9, -10, 26, -20, -27, -34, -46, 5, 2, -36, 1, -28, 7, 15, -3, 2, -23, 8, -1, 74, 6, 13, 15, -5, 0, -17, -5, 1, -4, -4, 4, -15, -11, -19, -17, -26, -5, -12, -16, -20, -26, -2, -12, 19, 6, 20, 0, 23, -20, -8, 10, 3, 15, 14, 15, 6, -1, -13, -26, -52, 15, 8, -14, 2, -3, -21, -18, -13, 11, 25, 8, 13, -4, 16, 10, 6, -6, -6, -8, 15, 11, -4, -8, -12, -13, -6, -6, -7, -46, -27, -6, 5, -12, 15, -6, -33, -10, 17, 1, -12, 24, 5, 15, -9, 5, -5, 6, -11, -3, 16, 10, -6, 3, -4, -26, -22, -18, -46, -11, 9, 4, 13, -10, -20, -27, 4, 10, 17, 12, -14, -3, 6, 46, -3, 18, -1, -13, 13, -14, 10, 7, -36, -3, 3, -62, -32, -6, -2, 2, 17, 1, -13, 6, -6, -2, 11, 0, 7, 33, 24, 21, 11, 38, -3, 18, 15, -2, -18, 11, -14, -15, -20, -12, -72, -30, 5, 23, 38, 17, -8, 7, 2, 9, 6, 20, 35, -1, 18, -19, 2, 53, 18, -2, -16, -7, -13, 9, 28, -5, -2, -6, -39, -28, -2, 1, 14, 20, -7, 2, -1, -30, 16, 23, -2, 9, -17, -15, 7, 26, -3, -1, 15, -13, 1, 0, 32, 4, 46, 10, 2, -1, -34, -21, 25, -42, 11, -3, 26, -6, 13, 0, 7, 11, -12, -22, -27, 14, 7, -8, 11, -1, 14, -22, -3, 29, 17, 11, -19, -11, -21, -3, 18, 3, -9, -12, -17, 29, 12, 4, 6, 1, 19, -3, -37, 4, 3, -11, 13, 17, -20, -32, 6, 17, 48, 28, -16, 1, 4, 5, -3, 17, -31, -70, -31, 24, 6, -11, -16, 10, 40, 0, 12, 36, -3, 1, 5, -11, 5, 27, -11, 35, 22, 6, 6, -3, -3, 4, 5, -14, -51, -47, -41, 30, 7, 8, -5, 6, 28, 6, 37, 57, 8, 17, -21, -1, 14, 8, 5, -1, 13, -45, -30, 1, 27, 24, 22, -12, -32, -67, -84, 16, 20, -14, 2, 8, 30, 31, 32, 24, 17, -16, 19, 7, 31, 35, -16, 2, -14, -49, -1, 21, 1, 11, 43, -6, -74, -112, -120, -3, 61, 11, 27, 9, 15, 8, 12, 24, 18, -4, 18, -15, 75, 37, -18, -34, -57, -101, 21, 34, 13, -7, 20, -6, -88, -113, -89, -10, 73, 31, 40, 32, 40, 28, 26, 61, 16, -5, -13, 17, 30, 17, -33, -49, -77, -77, 10, 54, 31, 48, 36, -13, -55, -85, -131, -30, 54, 27, 26, 47, 35, 29, 33, 48, 8, -7, 8, -9, -45, -15, -5, -35, -91, -95, 7, 41, 19, 23, 48, -15, -88, -91, -90, 10, 71, 62, 26, 10, 29, 41, 59, 78, -8, 8, -11, 20, 0, -23, -51, -67, -92, -84, 36, 43, 14, 33, 28, -28, -89, -115, -80, -44, 26, 52, 29, 26, 49, 58, 67, 63, 20, -6, 13, -19, 1, -44, -71, -66, -81, -51, 55, 43, 3, 44, 14, -64, -92, -83, -134, -52, 38, 44, 13, 26, 23, 20, 36, 32, 4, -2, 7, 21, 10, -35, -11, -43, -105, -31, 23, 37, 1, 36, 41, -71, -83, -104, -117, -89, -1, 28, 25, 51, 52, 19, 21, 46, -8, 10, -5, -7, -26, 19, -9, -57, -57, -25, 39, 24, 44, 74, -8, -88, -98, -88, -90, -50, -24, 38, 29, 9, 63, 38, 22, 1, -9, -10, -13, -8, -18, -3, -5, -60, -68, -46, 41, 41, 66, 45, -24, -56, -70, -100, -79, -92, -21, 43, 58, 52, 64, 27, 12, 8, 0, -12, 1, -9, 10, 28, 15, -35, -47, -60, 14, 13, 28, 54, -14, -53, -79, -117, -78, -110, -18, 47, 33, 51, 32, 18, -14, 1, 18, 10, -15, 17, 12, 38, 47, 47, 28, -29, 24, 31, 48, 44, -37, -17, -74, -71, -50, -72, -39, 22, -5, 25, 41, 54, -6, -34),
  19 => (15, 4, -16, -8, 8, 3, 12, -5, 5, -6, -7, 15, 4, -16, 6, -18, -13, 7, 12, 5, -10, -16, -18, 5, 16, 6, -15, 0, -18, 9, 3, 18, -14, 14, 15, -17, -17, 7, 9, -5, 3, -15, 14, 14, 8, -18, 17, 13, -12, -4, 13, -4, 14, -16, 8, -13, -19, -4, -18, -5, -3, -5, 14, 8, -3, 2, -4, 13, 4, 3, 5, -15, 5, 1, -19, 6, 12, 13, 11, -10, -10, -16, -20, -8, 19, -7, 15, -2, 4, 15, -7, -12, 22, -23, -6, -13, 11, -20, -28, 1, 10, -34, -6, -1, -25, 15, -14, 14, -1, 13, 17, -21, 20, 14, 18, -7, 6, -5, -5, -14, 12, -22, -11, -10, -21, -67, -43, -13, 0, -21, -20, 3, -5, 11, 2, 18, -3, 13, -2, -2, 0, -1, -5, -20, 7, -5, 0, 0, -5, -35, -4, -3, -19, -63, -47, -25, -24, -15, -10, -23, -18, -12, -16, -8, -13, 19, 0, 0, 5, 4, -2, -10, 15, 3, -4, -23, -25, -32, -32, -17, -54, -78, -39, -23, 0, -27, -48, -24, -4, -7, 3, 8, -10, 5, -7, 18, -3, -8, -1, -12, -16, 6, 15, -12, -23, -36, -41, -77, -37, -59, -88, -80, -52, -60, -62, -27, -47, -26, -4, 0, 14, -21, 6, 15, 4, -7, 5, 20, -14, -8, -25, -24, -32, -68, -88, -66, -30, -42, -64, -98, -91, -31, -54, -4, -22, -28, -14, -27, -22, -4, 7, 12, -12, -12, 20, -1, 0, -18, 1, 11, -36, -88, -56, -71, -46, -29, -54, -66, -70, -64, -34, -30, -47, -24, -9, -2, -24, 13, -20, 14, -3, 2, -6, -18, -15, 12, 6, -19, -34, -56, -35, -55, -39, -32, -53, -60, -27, -15, -40, 6, -47, -38, -34, -40, -2, 13, 7, 15, -13, -3, -17, 20, 19, 17, 0, 1, 2, 14, -6, -43, 12, 4, -41, -43, -33, -50, -40, 0, -6, -56, -52, 28, 2, -12, -11, 12, 4, 14, -18, 18, -16, 16, 21, -22, 9, -4, 17, 8, 6, 35, -4, 12, -22, 2, 9, 7, 5, -6, 10, 20, 28, 13, -19, -12, -10, -2, 11, -8, 17, -6, 15, -6, 11, 22, -12, 4, 5, -12, 24, -5, 0, -8, -3, 35, 19, -14, 9, 4, 11, 18, 3, 4, 10, -17, 13, 19, -10, 13, 20, 20, 21, 17, 17, -9, -12, 9, 14, -3, -21, -29, -29, -12, -12, -45, -35, 5, 4, -8, -14, -13, 0, 16, -19, -8, -16, 31, 21, 35, 16, 12, -4, -2, -27, 11, -14, -53, -37, -76, -64, -30, -30, -58, -27, -32, -2, 15, -6, -2, -1, -4, 9, 8, -24, 2, -12, 4, 5, 53, 19, 42, 25, 37, 28, -1, -5, -18, -22, -48, -43, -25, -15, -1, 4, -1, -20, 10, -10, -13, 3, -7, -25, 21, -1, 10, 19, 50, 60, 64, 39, 63, 36, 27, 7, -8, -9, 7, 2, 8, 23, 56, 49, 14, -6, -33, 14, 10, 8, 9, 13, 37, 32, 31, 4, 6, 13, 45, 48, 51, 10, 20, 1, -16, -3, -37, -13, 26, -5, 33, 39, 13, 16, 13, -14, 20, 4, -6, 0, -3, 25, -1, -4, 18, -1, 42, 51, 59, 18, 31, 11, 13, 11, -1, -1, -38, 0, -7, 4, 24, 30, 16, 2, 11, -4, 0, -22, -54, 5, -2, -10, 13, -10, 12, 4, 13, -7, 6, -5, 20, 11, 30, 21, -14, -27, -32, -15, -18, 21, 16, 0, -7, -10, -15, 5, -33, -58, -24, -68, -41, -21, -63, -54, -12, -13, -3, -11, 7, -3, -17, 22, 22, -17, -47, -21, 4, 26, 14, -11, -19, 18, -5, -42, -53, -1, 9, 11, 14, -21, -17, -14, -11, 15, -41, -35, -36, -13, -39, -6, 7, -16, -61, -40, -47, 8, 40, -3, 6, 20, -7, -34, -67, -17, 17, 2, 10, 17, -11, 43, -8, -13, 8, -9, 16, 14, -9, -20, -3, -14, -39, -24, -33, 23, 31, -21, -15, 17, 1, -7, -57, -12, -50, -7, -11, -20, 15, 17, 19, 11, -11, 6, 9, 11, -4, -34, 4, 30, 2, -31, -12, -29, 5, 4, 6, -4, 12, -24, -6, -7, -10, -13, -24, -1, -5, 37, 18, 14, -32, -24, -24, 9, 2, -14, -24, 24, -5, -26, -10, -24, 0, 18, 2, -17, 16, -18, -8, -7, -51, -16, -17, -16, 27, 6, 20, 4, 10, -17, -29, -23, -6, 14, -1, 19, 2, 7, -7, 0, -18, 20, -17, -3, -16, -1, 9, 1, -4, 24, -7, -9, 5, -19, 25, 9, -16, 2, 13, -18, -9, 5, -24, 9, 8, 13, -24, -14, -34),
  20 => (-5, 6, 16, 15, -6, -6, 9, 4, -7, -20, 5, -7, 19, 19, 11, -28, -36, -13, 29, 26, -10, 11, -4, 11, -20, 10, -4, 18, 1, 5, -4, -2, -20, -8, -8, -20, 17, -11, -5, 15, 6, 28, -7, -15, -36, -34, -5, -8, -39, -35, -37, 46, 43, 7, 1, 16, -13, 14, 2, -12, -7, -14, -11, 15, 1, -5, 23, 10, 11, -6, -40, -7, 3, 53, 6, -31, -23, -47, 32, 74, 48, 16, -8, 17, -12, -11, 6, 14, 20, -14, 4, -11, 8, -11, -20, 27, -9, -45, 2, -36, -6, 8, -57, -43, 6, -2, -15, 35, 79, 20, -18, -2, -17, 9, 20, 7, 16, -6, 9, -2, -7, -23, 0, -37, -67, -60, -32, -19, -13, -28, -9, 9, 18, 8, -2, -7, 2, 1, 4, 1, -5, -13, -2, 7, -6, -20, -18, -21, -36, -35, -32, -49, -73, -4, 16, 4, -40, -43, 31, 6, -5, -5, -30, -22, -35, -5, 3, 10, -2, -19, 0, -20, -4, -3, -1, -24, -32, -68, -49, -50, -20, 49, -25, -29, 13, -10, -14, -3, -30, -31, -2, -40, -44, -6, 2, -11, -7, 20, 9, -2, 16, 9, -14, -34, -35, -5, -53, -15, 67, 30, -14, -28, 19, -14, -39, -38, -19, -33, -34, -26, 21, -5, 74, 14, -1, 6, 1, 18, -1, 4, -24, -57, -18, -66, -61, 58, 66, 23, -10, 45, -7, -41, -33, -6, 30, 7, 31, -15, 11, 5, 64, 42, -1, -5, 18, -2, -15, 15, -9, -21, -32, -90, 27, 40, 27, 10, -14, 1, 11, -13, -37, 41, 72, 49, -5, 31, 0, 43, 33, 24, -10, -12, -4, 19, 4, 30, -14, -34, -81, -46, -15, 39, 86, 76, 10, -26, 11, -32, -55, 15, 25, 6, -5, 31, 37, 59, 43, 37, -17, 10, -12, -5, -3, 5, -63, 0, -51, 10, 32, 48, 78, 17, 9, -37, -22, -47, -12, 9, 21, 16, 40, 17, 52, 70, 63, 33, -5, -12, 7, 10, 16, 58, -21, -35, -45, 17, 25, 78, 67, 5, -21, -38, -30, -23, -22, 8, 36, 53, 59, 45, 47, 61, 59, 41, -14, 15, -8, 21, -6, 15, -42, -93, -9, 38, 46, 48, 27, -51, -62, -80, -5, 9, -13, 2, -1, 9, 45, 22, 48, 88, 45, 28, -4, 2, -8, -8, -9, 20, -71, -48, 13, 25, 27, 69, -2, -16, -40, -42, 36, 25, -22, 6, -11, -5, -22, -27, -3, 47, -13, -39, 15, -12, -4, 10, -9, -25, -80, -39, 22, 19, 43, 9, -4, -27, -22, -7, 10, 9, -10, 49, 14, -11, -14, -39, 2, 6, -3, -39, -20, 8, 0, 17, -58, -81, -127, -57, 6, 26, 32, -16, -31, -28, -51, -23, 13, -24, -19, 12, 17, -3, -2, -29, -7, 18, 22, -28, -7, -13, -14, 5, -42, -82, -114, -4, 56, 11, -3, -17, -22, -47, -41, 8, -7, 6, 4, 22, 11, -8, -9, -27, -28, -27, -13, -46, -6, 2, -5, -8, -33, -88, -96, 4, 36, 3, 12, -11, -11, -11, 14, 17, -1, 1, -10, 1, -10, -9, -36, -32, -59, -39, -20, -40, 3, 11, -9, -4, -9, -92, -79, -6, -8, -4, -15, 3, 6, -2, 2, 23, 19, -26, -26, -39, -46, -1, -37, -46, -16, -49, -69, -20, -19, 15, 20, 13, -13, -57, -30, 26, -28, -29, 16, 2, -1, 10, -2, 9, -15, 0, -55, -62, -54, -35, -55, -11, -85, -51, -46, -73, 3, -3, 12, -15, -18, 6, 8, -11, 14, -5, 25, -3, -24, -24, 0, 4, -38, -35, -66, -82, -84, -53, -43, -9, -7, -54, -31, -10, 10, -13, -11, -19, -47, -29, 14, 28, 11, -3, 43, -14, -7, -18, 5, -16, -57, -64, -93, -69, -83, -74, -76, -55, -22, -15, -30, -16, 8, 20, 20, -17, -30, -41, 3, -11, -4, 29, 11, 34, 17, 41, -4, 0, -52, -76, -78, -92, -62, -88, -63, -42, -22, 0, -9, -44, 10, -7, 3, -17, -45, -66, -1, 2, -29, 0, 1, 22, 26, 29, 12, -7, -30, -59, -81, -54, -25, -48, -67, -35, 5, -17, -11, -7, 1, -10, -10, -7, -3, -27, -29, -32, 16, 15, 46, 25, 25, 40, 16, -16, -12, -46, -31, -53, -44, -22, -53, -40, -22, -11, 13, 1, -10, -3, -11, 1, 20, -40, 5, -81, -10, 11, 37, -9, 9, 10, -19, -16, -22, -14, -61, -59, -27, -31, -1, 6, -16, -4, 27, 23, -13, 0, 2, 10, 20, -8, -13, -36, -11, 1, -3, -13, -33, -15, -31, -60, -73, -50, -74, -61, -12, -17, 12, 9, -10, 22, -13, 9),
  21 => (4, -3, 17, -14, -20, 9, -15, 6, -8, 5, 15, -13, 13, 18, 3, -34, -4, -33, -4, 23, 19, 10, -36, -20, 5, -10, -14, 5, 15, -16, 18, 10, 19, 12, 5, -1, -16, -16, -12, -2, 10, -29, -16, -62, -2, -26, 8, 14, -34, -28, -17, -8, -12, -19, 18, 11, -19, -8, -1, 20, 14, 1, -14, 1, -1, -9, 6, -21, -15, -63, -19, -32, -23, -22, 33, -11, -23, -17, 22, 37, 53, 17, -6, 14, -16, -5, 11, 16, -11, 6, 11, -2, 7, 10, -42, -30, -49, -43, -15, 1, -35, -71, -3, -16, -4, 1, 9, 36, 3, -6, 14, -16, 17, -16, 9, -20, -1, -17, -19, -17, 4, 40, 9, 6, -17, -28, 4, 8, 20, -7, 6, 27, 6, 11, 30, 75, 46, 16, -10, -1, -10, 12, -11, 19, -16, 12, -3, 9, -8, 35, 56, 43, 62, 48, 25, 19, -7, 29, 13, 36, 18, 31, 49, 79, 44, -38, -19, 0, -11, -13, -9, -14, 1, 12, -17, -16, 6, 48, 76, 51, 35, 45, 36, 28, 36, 25, 37, 40, 33, 14, 28, 22, 31, -9, 0, -4, -9, 1, 7, 10, -12, -1, -14, -45, 5, 7, 18, 24, -17, -11, 2, 32, 30, 21, 30, 31, 7, 12, -13, -1, 3, -20, 11, -13, -7, 16, -12, 9, -17, 20, -35, -50, -11, -77, -51, -77, -53, -62, -54, -28, -29, -47, -56, -64, -30, -26, -33, -75, -83, -30, -69, -22, 13, 6, -9, -13, -14, 7, -23, -33, -47, -63, -87, -64, -54, -29, -64, -67, -23, -56, -22, -44, -56, -62, -82, -106, -106, -53, -43, -29, 7, 6, 1, 6, -20, 6, -33, -21, -35, -21, -16, -36, -9, 0, 19, -19, -11, -6, -17, -14, -22, -39, -81, -75, -88, -59, -74, -55, -10, -18, 10, 0, -16, -49, -1, 42, 9, 30, 40, 44, 42, 53, 48, 26, 25, 3, -3, -27, -15, -57, -44, -21, -58, -40, -62, -32, 12, -8, -7, -13, 5, 31, 5, 1, -15, -16, 1, 10, 37, 5, 15, 31, 73, 54, 30, 31, 26, -21, 0, 14, -4, 0, -21, 9, 20, 18, -19, 15, 16, 15, 23, -35, -9, -27, -28, -30, -38, -28, -38, -9, -6, 34, 39, 33, 30, 2, 18, 51, 44, 37, 21, -29, 3, -12, 13, 19, 32, -26, 17, -12, 9, -18, -30, -24, -35, -61, -71, -53, -84, -62, -50, -42, -12, -6, 15, 23, 34, -4, 40, -27, 8, -7, -5, -15, 6, -48, 0, -21, -14, -14, -12, -33, -22, -1, -14, -45, -48, -69, -79, -58, -50, -16, -20, -6, 32, 49, 46, -13, -3, 1, 7, 15, -47, -77, 4, -12, -2, -26, -22, 27, 27, 24, 3, 16, 2, 2, 1, -6, -20, -19, -18, -37, 3, 30, 66, 22, 16, 1, 3, 14, -35, -67, -5, -21, 10, -22, 14, 2, 25, 22, 9, 21, 21, 35, 1, 26, 15, -16, -34, -21, -47, 29, 25, -22, -13, 18, -12, 15, -35, -52, -20, -21, 4, 16, 20, 3, -21, -24, -4, -8, -6, 9, 18, -5, -11, 33, 12, -8, -16, -19, -4, -41, -16, 14, 6, 11, -6, -31, -20, -20, 5, 13, 11, 0, -17, 0, -7, 3, -19, -6, 17, -19, 14, 24, 68, -9, -30, -62, -40, -46, -14, 8, 15, 11, -44, -4, -71, -24, -15, -17, -28, -53, -36, -30, -61, -30, -21, -40, 5, -1, -10, 6, 18, 15, -28, -58, -31, -18, -19, 17, -3, 17, 12, -35, -34, -36, -43, -34, -54, -45, -30, -26, -38, -50, -43, -35, -41, -10, -43, -18, 27, 26, 13, -28, -25, 16, -13, -1, 11, 8, 0, -44, -39, -36, -31, -11, -62, -75, -27, -30, -35, -17, -24, -12, -27, -16, -22, 2, 28, 28, 26, 32, -52, -13, 6, 3, 7, -6, -28, -12, 12, 22, 42, 17, 11, 16, 12, 17, 10, -3, 6, -11, -1, 7, -25, -9, -2, 2, 33, 10, -54, -26, 11, -10, 14, 1, -5, -5, 57, 51, 62, 19, 67, 51, 10, -1, 35, 25, -7, -2, 17, 9, 14, 24, -4, 25, -2, -41, -32, -57, 15, 17, -3, 3, 9, 30, 52, 65, 40, 42, 46, 23, 2, 22, 11, 18, 30, 16, 39, 43, 8, 23, 3, 11, -16, -18, -54, -56, -16, 7, 14, 0, 9, 9, 55, -2, 58, -14, -15, 13, 5, 5, 37, 48, 41, 73, 25, 54, 34, -19, -6, 31, 10, -23, -76, -45, 2, -13, 19, -9, -14, -10, 7, 2, -11, -10, 6, -14, -13, 22, 1, -21, 6, 0, -6, 9, 14, -46, -50, 9, 11, 11, -52, -21),
  22 => (-20, 15, -6, 10, 18, 10, -19, -13, 13, 17, -9, 16, 2, -7, -29, 15, 5, -21, -44, -52, -53, -6, -2, -4, 2, 14, -12, -13, -9, -7, -15, 14, -11, -18, -18, -9, -16, 6, 6, 1, -17, 52, 29, 27, -13, -16, -26, -62, 5, -13, -18, 50, -5, 2, 0, -20, -13, 16, -14, 19, -6, 15, 6, 19, 21, 3, -10, 25, 22, 18, -2, 9, 52, 43, 40, 27, 48, 39, 85, 71, 17, -20, 4, 18, -5, 19, -3, 15, -14, 1, 12, 8, -25, -10, 31, 28, 19, 3, 31, 13, 52, 32, 39, 43, 24, 48, 63, 68, 64, 56, 12, 11, -12, 3, -8, 4, 1, 2, 3, -9, -1, 64, 36, 40, 44, 37, 9, -13, 29, 27, 31, 23, -1, 34, 25, 35, 34, 22, -18, 10, -14, 8, 10, 11, -14, 2, -1, -2, -4, -6, 14, 40, 19, 7, 16, 2, 13, 33, 31, 27, 6, 10, 13, -10, -7, -10, 1, -18, -20, -10, 10, 1, 19, 11, 9, -20, 10, -2, 3, -3, -8, 8, 41, 42, 26, 57, 33, -27, -20, 0, -26, -37, -37, -2, 10, -16, -2, 1, 4, -18, -4, -19, 2, -7, 39, -19, -28, -22, -56, -34, -64, -77, -51, -49, -75, -97, -75, -76, -61, -93, -47, -21, -71, -38, -4, -5, 17, 8, -1, -18, -6, 39, 34, -30, 49, -1, -9, -8, -31, 7, 9, -35, -61, -59, -33, -42, -64, -95, -44, -43, -47, -32, 11, -2, 11, 6, 7, -3, 16, -7, 24, 21, 78, 25, 34, 22, 0, 35, 46, 35, -13, 18, -12, 2, -22, 0, -12, -21, -81, -44, -20, -11, -10, 2, 13, -27, 5, 1, 42, 28, 58, 30, 9, 11, -1, 10, 24, -6, -9, 14, 10, 9, 38, 39, 2, -5, -30, -27, 18, 0, -6, -15, 10, -64, -29, -24, -66, -24, -8, 1, 15, 32, 54, 46, 27, 15, 0, 29, 16, -3, 25, 22, 37, 12, -2, -6, 16, -1, 13, 6, -2, -18, -35, -24, -43, -43, -43, -54, -53, -33, 2, -12, 20, 19, 37, 75, 10, 2, 18, -7, 29, -23, 20, 18, 15, 8, 7, -18, -2, -44, -93, -60, -34, -9, -35, -49, -40, -85, -45, -32, -16, -24, -25, -3, 13, 2, -35, -37, -16, -37, -3, -17, 12, -5, 19, -20, -7, -36, -13, -39, -17, -28, -67, -77, -46, -75, -53, -37, -88, -62, -16, -1, 1, 1, -32, -48, -12, -41, 0, 5, 16, 10, 12, -6, -32, -28, -52, -30, -15, 13, -43, -20, -12, 3, -9, -31, -33, -50, -25, -23, -29, -32, -47, -3, -23, -30, -1, -16, 2, -15, -11, -18, -20, -38, -40, -36, -21, 5, 6, 25, 6, 29, 32, 0, -16, -23, -39, -3, 5, 2, 0, -25, -22, -23, 12, 12, 13, 17, -10, -4, -12, -45, -16, -43, -14, -14, 6, 29, 58, 11, 15, 25, -1, 28, 18, 5, 15, 16, -2, -20, -9, -11, -11, 5, -7, -16, 8, 18, 4, -30, -43, -27, -26, -9, 30, 66, 41, 27, 29, 2, 23, 55, 41, 18, -13, -2, -46, -41, -4, -4, -62, -22, -1, 16, 16, -11, 36, -55, -30, -24, -10, 1, 7, 18, 27, 25, 7, 2, 5, 42, 16, 4, 22, -25, -29, -36, -31, -2, -20, -27, -14, -12, 0, 20, -21, -24, -18, -27, -4, 12, 43, 16, 18, 19, 0, -38, -7, 0, -31, -20, -19, -22, -25, -21, -38, -26, 24, 14, -5, 11, -9, -18, -24, -45, -21, 3, 3, -11, 5, 2, 22, 15, -22, -40, -6, 39, 3, 9, -26, -26, -59, -53, -25, -3, 31, 55, 9, 16, -9, -3, -18, -29, -35, -27, -8, 12, 21, 39, 3, -9, -30, -67, 26, 57, 0, 12, -7, -25, -38, -63, 4, -7, 19, 7, -1, -14, 15, 2, -4, -57, -6, -7, 22, 34, 45, 33, 10, 30, -31, -60, 9, 40, 1, 24, -14, -46, -33, -31, -8, 13, 30, 1, -4, -10, 4, 8, 2, -8, 16, -4, -17, -5, 8, -14, 24, 42, -38, -38, 15, 19, -14, -6, 5, -22, -6, -27, 1, 2, -17, -33, 11, 12, -18, -8, 6, -9, -30, 15, 9, 18, 4, 21, -6, -12, -93, -27, -9, 12, 16, 4, -6, -35, -4, -23, 48, 4, -29, -28, 8, 14, -16, -10, -12, 1, 18, -19, -4, 27, 17, 40, -23, -57, -63, -76, 6, 25, 20, -8, 5, 22, 15, -3, 33, 24, -30, -11, -1, 10, 4, 4, 11, 16, 16, -24, -22, 1, 8, -23, 21, 28, 7, -23, 33, 31, 35, 7, 38, 58, 34, 48, 13, 16, -26, -14),
  23 => (7, 3, -6, -14, -2, -7, 17, -7, 0, 10, 2, -20, -13, -4, 17, -6, 18, 49, 26, 31, 8, -23, 3, 15, 21, 6, 0, 9, 5, 18, -5, -20, -9, 9, -4, 20, 19, 20, -17, -5, -9, -24, -42, 4, 13, 15, -1, -11, -42, -13, -20, -20, 10, -14, 11, -8, -19, 16, -4, -16, 8, 20, 20, -8, -19, 15, 8, -37, -53, -13, -16, -17, -53, -10, -13, -13, -8, -7, 8, 55, 21, 13, 5, -8, 12, -16, 4, -20, 2, 17, -16, 12, -7, -4, 7, -26, -15, -18, -2, -16, -31, -30, -50, -49, -9, -6, -13, 40, 48, 22, 7, -5, 20, -3, -9, -2, -17, -15, 4, 10, -10, -11, -22, -26, 2, -6, 26, 35, 37, -17, -18, -29, -6, 10, 22, 48, 86, 2, 1, 5, -2, -6, -19, 11, -17, 5, -18, -7, 14, -10, 35, 25, 34, 17, 29, 26, 43, 14, 10, -7, -3, 7, 22, 50, 61, 32, -13, -5, -6, -1, -3, 13, -12, 6, 12, 1, -24, 43, 40, 39, 33, -4, 13, 26, 30, -2, -5, -6, 14, 26, -3, 41, 52, 20, -32, 20, -14, -9, 7, 14, 12, 9, 12, -6, -34, 51, 43, 3, 10, -5, -9, 6, 14, 14, -8, 13, 2, -3, -35, 8, 30, -23, -15, 21, 7, -18, 11, 12, 11, 11, 25, -23, -7, 6, -14, -36, -29, -7, 33, 35, 32, 14, -18, 11, 46, 12, -12, -35, -59, -45, -30, 18, -1, 1, -3, -15, -1, -9, -8, -11, -27, -44, -50, -52, -35, -17, -19, 17, 31, 13, 2, 0, -5, 20, 10, -27, -31, -30, -43, 1, 20, -12, 18, -16, 2, -14, -9, -30, -56, -47, -100, -75, -1, -22, 6, -10, 16, -18, -14, -7, -14, 14, 43, -5, 14, -3, -46, -47, 11, 17, -17, -20, -11, -38, -15, -51, -65, -24, -16, -14, 2, 18, 6, 16, -20, -11, -10, 10, 9, 6, 39, -1, -16, -23, -27, -30, 6, -19, -7, -17, -17, -34, -13, -41, -30, -6, 9, 3, 12, 31, 6, 12, -14, -34, -12, 22, 1, 18, 20, -32, -54, -40, -8, -14, -17, 8, 20, -1, -19, -48, 15, -24, -5, 34, 14, 27, 56, 23, 27, -1, -17, 11, 32, 34, 31, 13, 15, -43, -31, -31, -45, -22, 16, 3, 1, -8, 4, -3, -13, -46, -23, -14, -25, 26, 20, -19, -27, 3, -17, -8, 26, 37, 9, 5, -2, -29, -45, 6, -12, -17, 8, -12, 3, 18, 21, 36, -7, -8, -15, -3, -34, -32, -29, -58, -30, -97, -74, -56, -19, 37, 15, -1, -2, -17, -24, -1, 7, 30, -4, 19, 20, 19, 48, 41, -8, -14, 30, -27, -17, -27, -45, -4, -41, -79, -73, -46, 9, 19, 19, -26, 20, -13, -54, -16, -36, 18, -15, -11, 7, -10, -1, -19, -47, -22, -11, -44, -15, -17, -15, -5, -19, -59, -35, -34, 40, 46, -11, -31, 55, 32, -27, -32, -18, -27, 8, -14, -6, 3, 49, 20, -30, -28, -40, -31, -20, -10, -25, -41, -43, -74, -91, -44, 19, 37, 47, 10, 40, 0, 20, -15, -24, -18, -16, 8, 8, -18, -39, -29, -31, -23, -52, 15, 14, 11, -44, -25, -39, -66, -103, -71, -36, 44, 66, 34, 13, 5, -18, -2, -2, 35, -6, -16, 1, 2, -7, -16, 30, -7, -18, 15, 40, 12, 14, 11, -41, -43, -82, -61, -10, 36, 66, 45, 50, 32, -53, -27, -12, 8, -5, -20, 3, 9, 15, -4, 14, 7, 22, 46, 40, 1, -10, -26, -35, -30, -37, -49, 6, 33, 57, 87, 71, 50, -1, -41, -32, 13, 3, -18, 12, -16, 0, 2, 31, 23, -9, -10, -10, 14, -6, -46, -43, -50, -66, -47, -30, 20, 70, 79, 67, 46, 3, -20, -8, 1, 9, 14, -10, 11, 29, 15, -14, -17, -18, 15, -13, -10, 37, 7, -15, 16, -42, -35, -10, 12, 29, 59, 45, 70, 8, -1, 23, 33, -6, 7, 7, 9, 8, -4, -8, -5, -23, -12, -31, -38, 21, 20, 8, 14, -8, -35, -53, -7, 24, 49, 56, 63, 33, 48, 12, 48, -9, 3, 17, 19, 19, -12, 5, -17, 5, -6, -60, -69, -11, -32, -17, -37, -34, -35, -6, 1, 43, 95, 75, 47, 82, 49, 9, 5, -5, -10, -3, -15, -19, -3, -18, -1, -2, -22, -15, 2, -29, -13, -36, -61, -70, -78, -32, 21, 50, 29, 59, 37, 53, 40, 48, 22, 19, 20, -3, 16, 16, -4, -17, -17, 1, -21, 0, -13, -42, -25, -38, -69, -69, -23, -51, -10, 38, 23, 24, 11, 24, 35, -7, -26),
  24 => (1, -18, 8, -3, 18, 18, 7, 7, 2, 17, 19, 3, 18, -6, -21, -1, 10, -11, -3, -7, -22, -22, 2, -16, 18, -6, -6, -17, -7, -18, 13, -2, -19, 4, -18, -3, 3, -20, 3, 15, 20, 13, -6, 10, -17, 17, 16, 29, 41, 24, 29, 4, -5, 13, -10, -10, -5, -20, -9, -7, -2, -18, -18, 2, -8, 0, 35, -16, 23, 10, -10, -22, -25, -25, -6, 42, 49, 74, 82, 16, 23, -3, -4, -16, -7, -20, 3, 2, -1, -6, 6, 2, 48, 15, 6, 11, 23, -12, -6, 4, 7, 10, 15, 32, 62, 61, 49, 26, -1, -4, -19, -20, 5, 5, 5, -16, -14, 7, 20, 22, 21, 89, 100, 86, -13, 15, -10, -19, 47, 26, 47, 30, -6, -38, -23, -42, -24, -9, -3, -14, -11, -3, -8, 8, 14, 4, 10, 1, 65, 84, 55, 20, -7, -5, -9, -6, 3, -22, -3, 4, -12, -30, -47, -87, -87, -6, -19, 2, -19, -2, -4, 15, -11, 12, 35, -29, 42, 56, 6, 21, 5, -8, -4, 3, 0, -13, -3, 4, -14, -12, -40, -60, -50, -44, -20, -11, -8, 20, -12, 5, -12, 13, 32, 9, 42, 34, 28, 13, 32, 11, -1, -3, 19, 24, 18, 17, 16, -12, -8, -29, -21, -54, -13, 11, -5, 14, 20, 15, 13, 9, 30, 29, 47, 18, 12, 2, 52, 28, 45, 18, 29, 14, 48, 42, -13, 21, 43, -9, 10, -10, 21, -8, -1, -16, 20, 10, 20, -17, -12, -27, 1, 3, -40, -21, -29, 1, 35, 23, 4, 22, 39, 29, 7, 13, 14, 1, 0, -13, -14, -13, 0, 0, -14, 1, -3, -28, -52, -78, -17, -45, -32, -40, -34, -59, -57, -38, -60, -51, -29, -43, -19, 4, 27, 2, 5, 12, -4, 12, 16, 7, 0, -6, -12, -67, -78, -45, -2, 47, 13, 14, -42, -27, -51, -77, -45, -70, -60, -99, -74, -82, -58, -50, -26, -27, -39, 2, -10, -18, 17, -13, 9, -56, -52, 8, -35, 0, 33, 39, 73, 47, 45, 41, 18, 5, -8, -81, -37, -46, -120, -67, -48, -51, -47, -4, -18, -16, -4, 20, -19, -15, -2, -13, -44, -17, -1, 4, 44, 58, 76, 81, 66, 34, 34, -2, -5, 17, -4, -57, -61, -75, -61, -48, 11, 0, 20, 20, -13, -8, -36, -22, -65, -37, -61, -68, -30, -8, 21, 39, 42, 50, 51, 33, -4, 10, 37, -22, -53, -88, -74, -30, -6, -5, 3, -16, -6, -20, -1, -5, -34, -34, -54, -51, -34, -75, -35, -14, -18, 26, 51, 27, 27, 18, 12, -8, 34, -5, -36, -64, 14, 19, 10, 18, 13, 22, 30, -4, 6, -35, -16, 14, -19, -28, -66, -82, -70, -51, -4, 14, 20, 21, 47, -12, 24, 28, -19, -40, -7, -17, -10, 20, 59, 54, 29, 19, 22, 26, 6, 34, 36, -7, -2, -43, -87, -28, -17, -11, 10, 23, 2, 0, 25, 32, 33, -40, 7, -12, -7, 4, 46, 32, 7, 23, 44, 18, 35, 15, 36, 26, 21, 12, -26, 13, 13, 3, -12, -2, 17, 14, 22, 42, 37, -2, 1, 12, -10, -1, 61, 5, -19, -10, -2, -19, 33, 2, 22, 23, 24, -9, 8, 7, 2, 4, 2, 31, -15, 0, -12, 34, 45, -24, -4, 4, 14, -4, 47, 49, -25, -30, -27, -18, -6, -25, 10, -1, -12, 7, 19, 12, 21, 5, 28, 44, 22, -13, 9, 28, 41, -56, 14, 15, -19, -16, 51, 15, -15, -15, -24, 3, -11, -24, 38, 17, -1, -12, -37, 3, 9, -4, -13, 12, 19, 28, 5, 30, 21, -39, -4, 13, 12, -1, 2, 1, -36, -56, -13, -31, -46, -50, 31, 15, 26, -4, 6, -1, -6, 4, -31, -7, 7, 29, 31, 31, 25, -14, 10, -10, 9, -16, -19, -53, -15, -35, 2, 20, -24, -38, -33, -33, -17, 2, 10, -19, -2, -4, -25, -22, 6, 24, 15, -17, -9, -12, -5, 17, -1, -6, 8, -35, 8, -5, 27, 16, 24, 14, -16, -26, -31, -40, -19, -42, -41, -48, -80, -62, -28, 13, -34, -26, -24, -29, 15, -21, 9, 11, -9, -34, 2, 9, -15, 24, 48, 37, 30, 28, 28, -31, -18, -21, -30, -46, -99, -91, -65, -24, 17, -41, -16, -59, 15, 19, -18, -12, -5, -2, -35, 6, -17, -15, 19, 8, 53, 35, 18, -8, -4, -24, 10, -36, -67, -79, -50, -8, -35, 11, -25, -27, -9, 20, 3, 17, -12, -16, -24, -25, -15, -15, 9, 37, 44, 25, 34, -18, 1, -2, -7, 13, -31, -7, -12, 3, -3, -39, -27, 3),
  25 => (-4, -2, 11, 0, -8, 16, 15, 0, -13, 4, -12, -5, -10, 0, 14, -22, -24, 1, 34, -3, -6, -21, -10, -13, 17, -6, 6, -11, 15, 7, -8, 1, -6, -7, 14, -3, 3, -4, -16, -18, -11, -45, -46, -33, -42, -37, -10, -7, -1, -28, 9, -7, 7, 0, -16, -16, -6, 9, 13, -17, -3, -16, 3, 3, -12, -25, -43, -41, -49, -7, 45, 29, -43, -51, -82, -41, -32, -49, -43, -45, -18, -17, -16, 2, 19, 2, -10, -20, 5, -14, 10, -9, -20, -31, -44, -4, 20, 58, 56, 15, -49, -35, -56, -12, -6, -51, -19, -38, 35, 11, 0, -1, 5, -10, 17, -9, -4, -6, 4, -2, -16, -74, -63, -8, 39, 25, 43, -9, -20, -32, -44, 2, -15, -33, -29, -11, 12, 34, -17, 8, -18, 16, -11, -14, -11, -11, -10, -25, -41, -33, 9, 15, 37, 9, -25, -32, -7, -14, -8, -5, -43, -53, -50, -1, 4, 3, -8, -11, 6, 1, 16, -1, 4, 6, -31, -21, 6, -24, -28, 38, 19, -62, -10, -8, 50, -3, 9, 17, -31, -76, -82, -30, 5, 31, -19, -8, -11, -7, -2, -19, -4, -19, -25, -37, -25, -64, -8, 19, -57, -37, -8, 17, 37, 5, 35, 26, -24, -85, -55, -18, 5, 87, -9, -20, 12, 10, 15, 9, -2, -12, -57, -45, -91, -37, -12, -45, -54, -21, -1, 11, 71, 40, 9, 18, -37, -32, -34, -42, 19, 63, 73, 7, -17, 19, 5, 21, 20, 12, -8, -43, -51, 18, 6, -53, -51, 25, -27, 29, 82, 31, 26, -4, -43, -31, -18, -17, 11, 86, 64, 18, -13, -16, -16, -18, -10, 50, 31, 8, 17, 75, 55, -11, -39, -37, -50, -40, 33, 56, 68, 36, -23, -1, 5, 23, 24, 37, 79, 34, -18, 20, 14, 20, -1, 27, 62, 47, 81, 50, 38, -15, -40, -25, -56, -41, 26, 67, 62, 43, 21, -5, -14, 21, 12, 36, 18, 13, -15, -9, 6, 6, 19, 5, 56, 59, 31, 26, 7, -16, 10, -18, -22, -3, -18, 82, 52, 36, 27, 13, -35, -30, -42, 10, 17, -2, 20, 15, -7, -18, 4, 18, 91, 46, 6, 29, 19, 4, 1, 17, -3, -22, 25, 68, 61, 55, 13, 20, 2, -41, -82, -1, 56, 28, 7, -13, 10, 13, -9, 35, 99, -8, -5, -1, 4, 8, 26, -9, -8, -42, -24, -5, 15, 20, -5, 9, 17, -24, -81, 4, 23, 44, 10, -11, -6, -16, -9, 51, 32, -25, 18, 41, 22, -19, -3, -20, -44, -94, -48, -41, -26, 40, 13, -17, -18, -31, -45, 22, 40, 21, 16, -4, 15, -3, -21, 57, 54, 21, 64, 51, 13, -8, 9, -21, -33, -99, -92, -60, -73, 15, 31, 8, -24, -9, -20, -19, -6, -3, -13, 5, -14, -10, -13, 39, 28, 10, 30, 40, 14, -14, -30, -7, -71, -108, -75, -52, -49, -1, 23, 13, 32, 18, -21, -27, 15, 7, 18, 3, 10, -6, -4, 21, 33, 14, 13, 6, 58, -6, 3, -22, -22, -50, -43, -60, -49, 18, 29, 53, 42, 0, 21, -17, 3, 17, -8, 2, 10, -8, 3, 14, 24, 25, 15, 36, 16, 12, -2, 29, 5, 14, -14, -52, -61, 6, -21, 34, 3, -9, -24, -40, -45, -26, -5, -5, -13, 14, -35, -45, -8, -9, 24, 25, 24, -11, -2, 30, 24, 33, 18, -47, -41, -35, -32, -22, -6, 12, -8, -27, -45, -22, 11, -15, -1, 5, -21, -23, -27, -90, -42, 10, -8, 23, 14, 32, 26, 21, 18, -28, -28, -13, -21, 5, -13, 27, -18, -32, -9, 30, 17, 12, 16, 20, -27, -22, -16, -34, -34, -22, -16, 0, -4, 49, 33, 29, 28, 14, -15, -17, 14, 11, -24, 26, 18, -32, -12, 22, -18, -12, 14, 18, -11, -9, -45, -67, -42, -57, -48, -54, -15, 38, 29, 31, 40, 45, 34, 31, 29, 34, 15, 26, 7, -7, -36, -28, -5, 11, -21, 18, 9, -43, -54, -78, -70, -40, -42, -77, 2, 8, 24, 0, 31, 38, 39, 28, 33, 0, 0, -19, 19, -29, -5, -11, -14, -7, -19, -8, -32, -9, -46, -70, -40, -53, -23, -59, -55, -17, -40, -16, -18, -2, -3, 0, -7, -10, 10, 29, 9, -5, -37, -22, 14, -9, -13, 5, 2, 15, -13, -25, -24, -20, -64, -47, -38, -57, -17, -46, 6, -13, 39, 35, 8, 5, 20, 14, 7, -6, 3, -23, -18, 3, -12, -3, -1, -20, -6, -22, -4, 2, 2, -65, -78, -81, -37, -28, -31, 4, 13, 9, 12, 12, 5, -4, -7, -22, 16, -30),
  26 => (2, 4, 17, -3, 17, -13, -12, 8, 1, -13, -9, -14, -1, -1, -3, 28, 20, 37, 11, 27, 42, 1, -16, -20, -16, 7, 20, 20, -21, 6, -8, -13, 5, -5, 20, -4, -16, -7, -13, -25, -28, -15, -51, 15, 67, 18, 72, 62, -9, -10, 13, 0, 1, 11, 0, -14, -2, -15, -11, 16, 16, 15, -6, -7, 2, 0, -10, -57, -10, -6, 38, 70, 44, 13, -10, 9, -41, -35, -44, 9, -21, 15, -11, -6, 2, -19, -1, 10, -11, -10, 15, -9, 13, -5, -19, 15, -7, 13, -1, 23, 12, -10, -1, -24, -17, -69, -61, -30, -5, 4, 13, 15, 19, 20, 13, -2, -19, 6, 17, -12, 20, 5, -18, -26, -37, -1, -14, 12, 8, -22, 5, -11, -26, -26, -61, -30, -24, -8, 5, -4, -9, 0, -20, 18, 8, 8, 13, -15, 11, 40, -3, -30, 17, -19, 12, 5, -5, -16, -9, 12, -20, -3, -46, -52, -7, 1, -5, -14, -10, -12, -10, -14, 12, -6, 16, -3, -2, 6, -2, 20, 10, -10, -12, -6, 27, 23, 3, 24, 7, 1, -48, -48, -40, -9, 4, -9, -1, -6, -13, -15, 6, 11, 16, 11, 0, 0, 36, 56, 38, 26, -20, 0, 30, 37, -16, 29, 59, 27, -25, -31, -57, 5, -2, 3, -11, -19, 6, -1, -5, 7, -18, -22, 13, 63, 68, 25, 11, -6, -6, -10, 37, 5, 26, 40, 9, -4, -35, -24, -25, -22, -10, 5, 3, 9, 18, -8, -20, 5, -3, -10, 10, 24, 15, -27, -8, 26, 61, 34, 36, 0, -2, 6, -1, -21, -39, -50, -35, -23, -16, -29, -3, -9, 7, 4, 19, 10, 2, -18, -5, -19, -32, -66, -28, 5, 57, 50, 33, 9, -1, 11, -9, -23, -32, -49, -16, -38, -14, -33, -6, -1, -7, -8, 15, -18, -46, -80, -65, -14, -34, -25, 16, 80, 53, 33, -4, -17, -4, 7, 6, -42, -28, -53, -28, -31, -35, -33, -11, 4, -3, 5, -9, -5, -54, -65, -64, -19, -17, -3, 5, 37, 34, 39, 9, -11, 10, -10, 44, 2, -31, -26, -24, 1, -27, -6, -12, -7, -9, -1, 10, -19, -33, -48, -44, -22, -39, 2, 11, -13, -34, 3, 13, -12, 16, 4, 6, 22, 2, -13, -27, -1, 33, 12, 0, 3, -11, 4, 18, -32, 0, -14, -64, -60, -29, -61, -97, -133, -101, -77, -48, -16, 11, 3, 8, 15, -17, 10, -51, -47, 3, -16, -7, 0, -11, 17, -12, -35, 26, 7, -70, -67, -76, -72, -95, -137, -116, -83, -40, -6, 23, 18, 11, 12, 3, 18, -57, -18, 13, -46, 7, 6, -11, -13, 11, 6, -17, -5, -42, -64, -49, 2, -10, -30, -27, -18, -28, 1, 13, 15, 35, 71, 40, -5, -34, -54, 23, -20, 19, -6, 10, 1, -31, -6, -14, 39, 14, 26, 79, 41, 33, 36, 27, 17, 7, 3, 12, -1, 37, 53, 67, 28, 1, -47, 3, -12, 17, -15, 19, 7, -12, 7, 31, 69, 30, 19, 34, 23, -7, 6, 4, 37, 2, 6, 4, -8, 22, 63, 23, 27, -8, -35, 0, -29, -1, 0, 12, -5, -37, 3, 44, 33, 20, 10, 0, 28, 24, 40, 34, 34, 39, -8, -23, -33, 2, 30, 13, 35, 1, -16, 14, -10, -9, -14, 16, 3, -33, -13, 27, -2, 6, -3, -12, -13, 34, 18, 13, 51, 39, -16, -18, -17, -30, 10, 33, 15, 19, -13, 19, -18, -1, -13, 15, -20, 10, 32, 34, 16, 14, 9, 45, 30, -6, -16, 21, 31, -4, 13, -22, -42, -60, -24, 14, -3, 4, 3, -6, -11, 3, -1, 9, 12, -6, 26, 27, 35, 54, 40, 16, -1, 0, -1, -33, 2, -3, -40, -21, -26, -50, -55, -5, 27, 57, 40, 15, 12, -2, -11, 7, -12, 0, -37, 4, 17, -17, -20, -73, -35, -38, -63, -62, -47, -67, -34, -91, -49, -88, -32, 8, 64, 48, 39, 34, 42, 1, 16, 13, 18, 4, 4, -17, 13, -29, -42, -48, -28, -48, -69, -77, -64, -67, -87, -58, -64, -50, -33, 18, 20, 53, 26, 11, 44, 19, 9, -3, -8, 15, 15, -2, -32, -23, -17, -36, -13, -44, -29, -22, -31, -45, -43, -25, -25, -16, -1, 11, 44, 55, 28, -2, 18, 10, 13, 12, -13, 2, -7, -6, 5, -31, 11, -40, -22, -39, -43, -37, 7, -14, 13, -16, -29, -35, -21, -17, 20, 50, -7, 18, 11, -14, 16, -16, -6, 17, 8, -9, 14, 12, -14, -23, -1, -40, -40, -29, 9, -2, 21, 43, -7, -26, -18, -12, -15, 15, 13, -13, 21),
  27 => (-16, -11, 0, -16, 9, 14, 20, 14, -20, -3, 17, 2, -8, -9, -38, 57, 48, -7, -33, -10, 9, 29, 37, 10, -16, 0, 0, -4, 8, 14, 1, -12, 4, 15, -12, -8, -5, -11, -10, 18, 38, 31, 52, 27, 22, -8, -16, -37, -15, -25, 13, 17, 38, 18, 15, -1, 19, 12, -12, 21, -9, 16, 19, 9, 0, 10, 13, 41, 24, 9, -12, 32, 45, 25, 14, 38, -8, 31, 60, 71, 46, 25, -5, 7, 3, -8, -13, 17, -11, -13, 2, -9, 10, 13, 61, 18, -5, 0, 3, -6, 31, 9, 14, 23, 39, 45, 71, 79, 27, -9, -10, 5, -17, -16, -2, -13, 2, 19, -9, 6, 16, 107, 43, 78, 30, -1, 24, 25, 17, 29, 30, 46, 36, 32, 19, 8, 54, -33, 6, 3, -3, -11, -15, -17, -17, -12, 0, -19, 22, 38, 58, 89, 81, 48, 30, 34, 43, 23, 13, 27, -21, -7, -16, -19, -3, 4, -19, 20, -17, -3, 8, 11, -20, -14, 24, -19, 0, 10, -4, -31, -7, -37, -71, -64, -50, -28, -39, -31, -59, -71, -97, -103, -30, -4, -8, -16, -10, 4, -8, -13, 3, 4, -2, 1, -4, -50, -83, -127, -97, -61, -41, -46, -14, -21, -14, -30, -33, -44, -74, -60, -50, -20, -19, -10, 3, 8, 15, 17, 9, -6, 7, 22, -21, -62, -37, -41, 25, 41, 22, 20, 25, 9, -11, 14, 5, -44, -16, -2, -5, -43, -33, -30, 21, 16, -14, -13, -7, -14, 12, 40, -9, 22, 21, 40, 19, 27, -2, 3, -6, -4, 19, 18, 1, -10, 2, 40, 27, -16, -52, -1, 8, 20, 4, -15, 1, 9, 49, -16, -4, 35, 47, 29, 25, 45, 8, 12, -14, -18, -5, 28, 4, 9, 26, 18, 46, 27, -4, -4, 5, 0, 8, -5, 17, 1, -17, -38, -22, -46, -22, -9, 1, 12, 21, 35, 53, 16, 54, 49, 20, 24, 7, 24, 32, 3, 2, -19, 0, 0, -9, 10, -35, -30, -11, -16, -11, -37, -32, -28, -67, -52, -72, -54, 26, -12, 34, 10, 1, -18, 26, -7, 9, -12, 14, 11, 16, -10, 6, 5, 0, 14, -13, -3, -8, -25, -15, -21, -35, -47, -33, -49, -71, -62, -44, -43, -35, -29, -30, -19, -31, -43, 8, 8, 17, 17, 3, -1, 7, -50, -86, -33, -65, -33, 14, -13, 8, 37, 25, 7, -14, -32, -13, -19, -43, -53, -46, -65, -30, -44, -7, -15, 6, 1, 3, -11, -6, -45, -71, -52, -26, -33, 21, 13, 8, 24, -2, -23, -25, -5, 34, -1, -7, -10, -18, -40, -22, -27, 11, -32, -12, 12, 16, 17, -15, -33, -56, -29, -46, -17, 4, 10, 17, -3, -37, -24, -15, -28, -14, 17, 5, -44, -3, -34, -28, -15, -16, -41, -20, 5, -2, 8, 23, 16, -21, -20, -31, -14, -31, -55, -27, -32, -9, -32, -22, 3, -12, 2, 3, 6, 45, 9, -9, -41, 2, -18, -21, -15, 4, -10, -14, 19, 20, 0, -33, -42, -62, -69, -66, -97, -35, -53, -12, -20, -7, 1, 18, 12, 21, -20, -8, -19, 14, -32, 3, 7, 1, 2, 27, 26, 1, -22, -17, -18, -93, -117, -113, -103, -111, -68, -3, -14, -19, 33, 32, 14, 8, 24, -15, -13, 29, -12, -13, -12, 12, -2, -29, 2, 18, 8, -36, 3, 10, -31, -22, 6, -4, 36, 63, 19, 4, 5, 30, -12, 20, 20, 7, 10, 42, 2, -9, -8, 19, 7, -30, -26, 34, 1, 22, 19, 51, 40, 37, 58, 71, 51, 47, 3, 11, 33, 49, 21, 23, -18, 11, 17, -19, 47, 4, 0, -8, -4, -31, -32, -8, 43, 41, 43, 33, 52, 24, 43, 12, 20, 5, 15, 21, 26, 52, 8, 48, -21, -11, 20, -16, 30, 2, -2, 19, 2, -17, -20, -3, -27, -5, 14, 44, 47, 37, -3, 20, 17, 16, 20, 11, 35, 16, -5, -3, -4, -42, -1, -13, 20, 6, -11, 7, 15, 7, -18, 0, 13, 29, -9, 2, 35, 21, 39, 24, 38, 36, 21, 36, 32, 39, 1, 2, 18, 7, -24, 15, 39, 17, 4, -14, -4, -9, 13, 28, 42, 9, -5, 1, -35, 24, 38, -11, 21, 44, 19, 52, 55, 48, 15, 14, -21, -2, 3, 29, 77, -20, -12, 11, 17, 18, -7, -20, -10, 13, -3, -10, -6, -20, -25, -49, -39, -41, -15, -5, 19, -5, -26, -21, 10, 42, -2, 34, 19, -10, 7, -11, 10, 7, -3, -12, 11, 10, -14, -52, -33, -78, -76, -56, -102, -42, -35, -23, -31, -33, 23, 29, 12, 52, 46, -2, 16),
  28 => (16, -4, -13, 8, -18, 11, -10, -2, 15, -6, 12, -11, 13, -17, -34, -17, -15, -7, 18, -12, -48, -18, -19, 19, 13, 7, 21, 9, 9, 3, 0, 6, -7, -7, -5, 18, -18, 17, -23, 11, -15, 10, 4, 12, -1, 19, 21, -14, -3, -11, 1, 4, -6, 15, -18, -10, -17, -6, 6, 2, 15, 17, 16, 1, 18, -17, -3, 25, -15, -38, -54, -24, 50, 78, 27, 3, 4, 6, 22, 11, 3, -14, 11, 3, 12, -6, -18, 2, 9, -19, -4, -14, -11, 0, 24, 28, 15, 10, 44, 17, 40, 30, 18, -36, -19, 7, 16, 17, -16, 17, 2, -6, 16, -15, -7, -1, 8, -10, -1, 3, 36, 14, -6, 2, -18, 47, 32, 37, 41, 5, -20, -32, -14, -1, 59, 40, -19, 9, 7, -3, 6, -9, -11, 13, -19, -5, 4, 39, 4, -49, -30, -28, -8, 13, 34, 4, 34, -26, -37, -69, -46, -4, 18, 13, 16, -6, -2, -6, -8, 15, -18, 2, -4, -16, -14, 29, -6, -9, -2, -24, 21, 12, 10, 6, 3, -8, -50, -58, -54, -7, 30, -14, -12, -23, -7, 8, -6, -3, 13, -2, -14, -14, 5, 40, -5, 4, 14, 1, 7, 31, 10, 3, 16, -22, 9, -61, -21, -15, -19, -21, -10, 5, -10, 5, 11, 4, -17, -2, 0, 7, 5, 21, 33, 33, 25, 12, 31, -11, 8, -6, -14, -32, 11, -61, -56, -66, -78, 6, -15, -11, -11, -7, 17, 18, -14, -13, 7, 6, -47, 16, 64, 40, 13, 16, -1, 1, -27, 2, 22, 5, 27, -46, -55, -41, -16, 16, -56, -3, -9, 16, -16, 4, -15, 10, 15, -4, -52, 21, 26, 38, 33, 19, 5, -22, -33, -20, 5, 8, 34, -28, -22, -15, -39, -7, 11, -28, -7, -14, 2, 19, -18, -16, -16, -36, -54, 1, -3, 38, 47, 35, 3, -49, -24, -61, -64, -35, 2, -50, -47, -33, -18, -16, -20, 3, 11, -3, -18, -4, 3, 6, -3, -79, -56, 35, 20, 17, 66, 38, -32, -56, -55, -35, -36, -49, -35, -2, -37, -33, -54, -1, 4, 17, 5, 18, 13, -20, 5, 15, 0, -112, -30, 13, 58, 65, 58, 65, -21, -55, -14, -47, -23, -14, 3, -7, -35, -33, -28, 2, 19, 0, 25, -4, -2, -18, 13, 10, -15, -94, -106, 39, 34, 22, 39, 24, 33, -35, -22, -24, -26, 3, 32, 8, -54, -55, -39, 8, 19, -5, -9, -17, -20, -8, 0, -3, -71, -120, -76, 18, 35, 15, 53, 38, -19, -35, -33, -28, -35, -21, 10, 0, -16, -33, 24, 15, 10, -24, -21, -9, 11, 0, 18, -13, -36, -143, -79, 22, 13, 42, 55, 48, -6, -45, -41, -26, -37, -52, 8, 13, 3, 2, 7, 27, -6, -33, -47, -27, 14, 19, 10, -9, -47, -142, -56, 15, 16, 56, 56, 45, 40, -33, -21, 1, -14, -14, 12, 27, 4, 1, -33, -48, -30, 2, -24, -20, 18, -10, 8, 20, -45, -119, -39, -9, 30, 35, 12, 36, 27, -53, -14, -13, -23, -26, 21, 32, 20, 5, 1, 10, -35, -1, -32, -17, 3, 16, 5, 3, -42, -114, -33, -1, 20, 24, 34, 36, 13, -23, 20, -24, -15, -17, 4, 2, 7, 12, 7, 8, 11, 2, 4, 11, -2, -3, -9, 0, 1, -76, -41, 8, 30, 31, 83, 69, -7, -14, -16, -22, -7, 1, -17, -3, -28, 28, -34, -34, 8, 24, 6, 25, -19, -19, 20, -10, -60, -51, -39, 0, 8, 10, 23, 31, -5, -31, -8, -2, -32, 5, -53, -10, -65, 9, 0, -15, -41, -2, -8, 16, 14, -2, -18, -13, 3, -16, -45, -17, 50, 31, 38, 8, -5, -24, -23, -18, 8, 21, -36, -81, -71, -30, 8, 10, -31, -3, -13, -13, 7, -19, 2, -15, -7, -28, -26, -42, -4, 44, 67, 48, 30, 8, -24, -4, 16, -12, -70, -102, -74, -47, -15, -7, 4, 3, -18, -4, -19, -4, 10, 1, -18, -1, 1, -33, -15, 52, 52, -8, 21, -10, 10, -1, -8, -37, -98, -80, -70, -29, 24, 2, -10, 16, 19, -15, -15, 19, -12, 0, -33, -9, 9, -26, 3, 27, 43, 34, 1, -32, -40, -38, -25, -43, -105, -54, -57, -37, -14, -23, 2, 19, -14, -16, -2, 0, 9, 4, -29, -3, -21, -71, -1, 17, 30, 5, 24, 7, -7, -31, -29, -45, -89, -52, -38, 1, -23, -12, -7, -9, 0, -17, 1, 17, -12, 13, 14, 1, 38, 25, 12, -16, 19, 29, -2, 28, -4, 2, -15, -40, -49, -6, 7, 9, -22, -10, -6, 16, 13, -7),
  29 => (5, -20, -8, 0, 8, 14, 20, 18, -6, 8, 7, 0, -20, -5, -19, 13, -47, -13, 29, -36, -44, -16, 11, -13, -8, -5, -18, -3, 7, 17, 6, -12, -11, 16, 10, -2, -15, 15, -14, -29, 3, -2, -17, 7, -22, -12, 2, -42, -35, -42, -44, 4, -5, 9, 11, 10, -9, -19, -9, 7, 9, 5, -13, -2, 11, 7, -13, 21, -17, -22, 4, 2, -8, -7, 8, 11, 11, 26, 13, 37, -1, 10, -13, -15, 3, 0, 0, 7, 1, 12, -8, 4, -22, -19, 46, 17, 11, 18, -31, -51, -50, 23, 6, 53, 12, 30, 22, -19, 2, 18, -20, -7, 16, 15, 7, -18, 4, -17, 17, 17, 1, 51, 49, 41, 50, 7, -4, -31, -36, 2, -23, 4, -6, 47, 31, -2, 15, -21, -13, 17, -19, -13, -17, -5, 16, 18, 27, -4, -20, 42, 18, -9, -7, -31, -37, -57, -42, -24, 15, -33, -3, 25, -1, -1, -10, -15, -1, 15, 4, -15, -13, 3, 15, -20, 18, 23, 1, 7, -14, -26, -25, 2, -34, -46, -37, -27, -15, -12, 2, -3, 7, 18, -71, 0, -6, 3, -12, 7, -1, -14, 5, -9, 5, 3, 35, -7, -18, -1, -20, -48, -46, -51, -34, -6, -18, 7, -12, -29, -17, 10, -41, -40, 1, 34, 14, 18, -15, 17, -5, -17, 42, 41, 18, 4, -5, -17, -20, -61, -75, -14, 16, 30, 28, -7, -17, 46, 35, 17, 7, -10, -11, -4, 11, 10, -19, 8, 8, -10, 15, 17, 13, 23, -21, -6, 4, -19, -6, 21, 10, 43, 46, 13, -1, 30, 3, -7, 33, 5, 43, 14, -1, -8, -18, -7, 17, 55, -5, -7, 11, 27, 13, 32, 30, 26, 39, 22, 46, 31, 9, 12, -6, 27, 24, -30, 21, -20, 31, -7, -7, 9, 2, -7, -10, 83, 9, 28, 32, 16, 37, 25, 22, 65, 49, 53, 50, 67, 45, -3, 19, 12, 9, -4, 13, 15, 12, 48, 6, 10, 5, 15, 19, 83, -14, -35, -53, -17, -17, -2, 24, 59, 52, 41, 37, 57, 22, 30, 28, 35, 25, -1, -3, 2, 25, 15, 17, -17, 11, -19, 31, 57, -38, -32, -64, -22, -1, -8, 40, 82, 71, 48, 46, 42, 28, 25, 6, 29, 42, 45, 16, 26, -16, -11, 1, 10, 7, -7, 57, 55, -33, -32, -27, 0, 25, 24, 75, 74, 44, 30, -15, 9, 0, 2, -39, 40, 14, 21, 18, -16, -14, -3, 0, -13, -11, 1, 29, 18, -4, 26, 13, 22, 51, 66, 58, 36, 33, 2, -11, -31, -12, -20, -39, -1, -3, -20, -28, -40, -5, -17, 10, -10, 2, 5, 37, 46, 13, -7, -11, 7, 20, 43, 44, 20, -10, -26, 19, -18, -38, -30, -41, -41, -10, -45, -38, -21, -20, -30, -18, -8, -8, 17, 17, 64, 29, 16, -15, 19, 18, 19, 22, 7, -21, -49, -37, 7, -36, 7, 11, -9, -56, -79, -49, 11, -42, -8, 8, 13, -20, 15, 15, 61, -19, 3, 31, 18, 49, 31, -12, -37, -30, -59, -39, 2, -14, -41, -5, -26, -39, -91, -86, -32, -52, -24, -10, -12, 17, 0, 48, 67, 10, 12, 45, 37, 8, -8, -4, -25, -12, -36, -43, -39, -30, -49, -24, -78, -71, -68, -34, -74, -27, 14, 19, 4, -14, 12, 44, 70, 12, 20, 26, 25, 30, 6, -25, -39, -42, -35, -56, -46, -78, -89, -59, -77, -96, -90, -74, -48, 0, 13, 10, -18, -10, 1, 17, 80, 7, 25, 32, 56, 37, 0, -65, -11, -24, -30, -41, -52, -66, -103, -59, -72, -62, -47, -53, -31, -41, 19, 14, 16, -11, -5, 55, 56, 14, 49, 18, 10, -14, -24, -54, -16, -15, -46, -51, -65, -76, -76, -35, -65, -68, -56, -30, -6, -12, -12, -10, 12, 1, -2, 37, 31, 44, 33, -5, -8, -50, -54, -40, -27, -44, -37, -55, -56, -55, -85, -67, -60, -61, -45, -13, 13, -18, -31, -14, -10, -11, -3, 34, 30, 38, 18, 1, -27, -42, -35, -41, -25, -58, -38, -64, -55, -55, -23, -39, -52, -66, -37, -26, -13, 17, 13, 12, 0, -11, 2, 17, 33, 33, -7, -7, -23, -20, -23, -57, -9, -10, -14, -44, -21, -60, -52, -50, -41, -14, 10, -15, 11, -8, 11, 17, -21, -20, -14, 3, 24, -8, 17, 7, -28, -30, -25, -25, -13, 15, -21, -57, -41, -42, -36, -36, -15, -22, -18, -14, 4, -10, 19, -20, -15, -13, -12, -4, 13, 18, 32, 3, -22, 17, -35, -18, -47, -39, 1, -37, -16, -23, -16, 3, 14, -7, 18, -11, -19, -8, -8),
  30 => (16, -16, 3, -7, -20, 6, -9, -18, 13, -20, -4, -19, -8, -10, 32, -19, -34, -65, -39, -38, -40, -4, 16, 14, -11, 7, -7, 12, -19, 16, 20, -6, 10, 0, 18, -8, -7, -17, 2, 29, 45, 31, 24, -7, -12, -22, 3, -3, -22, -8, 31, -5, 7, 8, 3, -12, -18, -8, -10, -11, 16, 19, 6, -20, 14, 44, 61, 38, 27, 22, 48, 40, 40, -5, 13, 4, -8, -31, -22, 8, 19, 16, 14, 9, 10, 17, -10, -12, 9, 5, -11, 16, 52, 67, 18, 25, 22, 32, 3, -9, 19, 7, 23, 16, -16, -17, -8, 7, 6, 3, 11, 18, -7, 19, -14, -20, 6, 3, -5, -8, 51, -11, 18, 7, 14, 39, 24, 18, -16, 27, -6, 9, -11, -40, -7, 5, -34, -55, 18, 1, 19, 4, 17, -5, 18, 17, -12, 52, 12, 8, 11, 6, 25, 14, 27, 2, -47, -16, -22, -11, -6, -35, -45, -9, -66, -9, -8, 18, -1, 15, 18, 14, -5, -17, 44, 81, 26, 22, 32, 46, 46, 39, 0, -25, -36, -22, -53, -20, -24, -46, -6, -33, 6, 2, -5, -14, 20, -9, 11, -13, 1, 2, 50, 75, 36, 35, 47, 18, 34, 2, 12, -4, 0, -10, -52, -13, 6, -5, -18, 21, 36, -17, -40, 5, 4, 16, -14, -8, 2, 3, 21, 58, 18, 31, 12, 6, 14, 1, 18, 32, 2, 5, -33, 0, -3, 25, 17, 13, 56, 8, -10, 11, -15, 0, -20, 13, 4, -2, 34, 9, 21, 0, 17, 21, -2, -8, -30, -18, -8, 4, 9, -16, 28, 55, 37, 34, 46, 33, -5, -12, -2, -15, 3, 7, 17, -17, 22, 3, -5, -8, -9, 6, 0, -8, 23, 42, 41, 38, 40, 23, 29, 51, 57, 42, 77, 41, -5, -27, 16, -17, 3, 11, -17, -9, 21, 10, -27, 12, 5, -17, 27, -16, 25, 38, 30, 33, -7, 55, 10, 69, 47, 45, 84, 33, 41, -9, 9, 4, 9, 0, 55, 21, 100, 31, 29, 25, -18, -15, 12, -3, 21, -1, 19, -2, -3, -2, 23, 14, 35, 29, 65, 60, 31, 7, 0, -10, -14, -12, 46, 39, 84, 51, 39, 51, 45, 23, 13, 19, 15, 14, 20, 45, 26, -5, 25, 31, 56, 52, 2, 78, -9, 15, -9, 17, 6, 4, 5, 37, 89, 86, 98, 31, 50, 56, 44, 52, 64, 58, 60, 63, 60, 32, 78, 42, 52, 12, 50, 31, 16, 22, 14, 7, 16, -6, 15, 44, 48, 80, 96, 39, 47, 58, 90, 83, 65, 75, 81, 82, 80, 86, 97, 69, 44, 23, -10, 2, -1, 4, 14, 16, 5, 18, 30, 33, 49, 69, 43, 38, 65, 43, 92, 80, 62, 36, 75, 32, 60, 41, 79, 74, 22, 2, -37, -15, -29, -13, -10, -15, 10, 21, 7, 37, 35, 53, 53, 23, 33, 17, 68, 54, 23, 33, 31, 59, 31, 26, 27, 49, 4, -11, 2, 3, -11, -12, 20, 18, -8, -4, 15, 7, 42, 35, 55, 3, 6, 11, 40, 40, 11, 30, 6, 40, 50, -2, 10, 0, -10, -4, -2, 3, 9, 16, 1, 11, -1, -2, -40, 12, 27, 32, 26, 4, 16, 28, 11, -2, 39, 6, 23, 16, 32, -10, 27, 16, -17, -22, -29, 1, -7, -7, 19, 17, 4, -1, -35, 5, 5, 19, 21, -14, -1, 39, 6, 15, 20, 28, 1, 19, 2, -7, 18, -5, 17, 9, -32, 2, -41, -5, 0, -4, -8, 15, -17, 6, 7, 14, 28, 21, 10, 1, 3, 10, 32, 29, 10, -6, 16, -13, -9, -40, 3, 5, 24, 7, 20, -1, 17, 3, -7, -19, 6, -5, 21, 25, 26, 6, -2, 22, 8, 3, 3, 3, 15, -13, 17, 1, -2, 2, -25, -33, -9, 9, -29, -40, -10, -1, 20, 1, -29, 1, 55, 53, 29, 37, 21, 6, 2, 38, -4, 18, 26, 7, -6, 10, 18, 17, -18, 7, 19, 2, 14, -39, 12, -11, -7, 4, 26, -6, -9, 32, 56, 25, 32, 15, 52, 29, 40, 32, 23, 32, -21, -1, 28, 28, -12, -29, 23, 9, 26, -51, 19, -7, 5, -15, -46, 12, 30, 6, 32, 4, 1, -3, -2, -24, 4, 1, 35, -2, -25, 3, 20, -17, -10, -8, 24, 30, 15, -40, 1, -21, 6, -20, 3, 64, 18, -45, -13, 34, -23, -12, -24, 2, 18, 22, 11, 13, 5, 3, 32, 4, 14, 11, 16, 3, 20, -16, -20, 10, 10, -11, -14, 45, 59, 43, 26, 13, 5, 26, -1, -16, 30, 58, 31, 39, 46, -12, 5, -16, -11, -40, -30, -20, -67, -35),
  31 => (2, 9, 11, 13, -12, -19, 19, -19, -3, 11, 8, -16, 21, 7, -1, -46, -28, -35, -13, -56, -48, -40, -25, 15, -8, 5, 3, -1, -2, 9, 2, 6, -20, 7, -3, -12, -6, -17, 8, 50, 50, 70, 45, 18, 4, 13, -17, -33, -18, -15, 15, 3, 24, -9, -20, 4, -4, 16, -13, 8, 1, -13, 17, -4, 11, 16, 93, 50, 47, 62, 28, 14, 16, 21, 10, 27, 18, 10, -35, -6, 0, -14, -7, -7, 2, 16, 19, -14, 19, -10, -19, -14, 36, 74, 89, 116, 106, 79, 37, 2, -30, 0, -3, 46, 34, -11, 8, -11, -2, -19, 14, 20, 6, 4, -15, 20, -17, 11, -4, 41, 83, 65, 96, 89, 76, 32, 15, -30, -26, -11, 19, 6, 19, -13, 25, -11, -23, -2, 5, -7, 5, -9, 13, -15, 2, 18, 31, 59, 49, 67, 53, 100, 51, 11, -8, -4, -19, -29, 1, 13, 23, 14, -19, 10, 4, 0, -2, -16, 8, 19, -18, 16, 10, -8, 34, 109, 53, 65, 82, 90, 42, 12, 13, 6, 9, -22, -21, -4, -11, 36, 40, -9, 15, -17, -11, -17, -5, 7, 15, -1, 19, -11, 80, 59, 81, 56, 35, 22, 38, 21, 18, -13, 2, -27, -41, -23, -12, 50, 0, 2, 1, 0, 11, -26, -10, 3, 8, 7, -20, -2, 56, 64, 55, 0, 17, 14, 34, 69, 51, 37, 17, -29, -9, -31, 2, 14, 17, 3, -8, 1, 4, -29, -15, 2, -20, -8, 19, -18, 39, -12, 6, -27, 4, 0, 28, 41, 31, 10, -9, -5, -13, -1, -7, 1, 17, 22, 1, 9, -3, -2, -17, -2, 7, -3, 11, -51, -13, -55, -54, -48, -24, -18, 48, 25, 17, 18, -10, 12, 0, -18, 14, 15, -6, -8, -38, 29, 3, 1, 16, 6, 16, 15, -9, -56, -66, -93, -107, -54, -24, 1, 16, 5, 24, 69, 49, 61, 13, 28, 45, 49, 20, -19, -59, -2, -12, 3, 8, 1, -3, 10, 0, -33, -35, -85, -70, -44, -20, 0, 9, 1, 40, 50, 47, 26, 52, 33, 62, 59, 24, 5, -57, -6, 32, 0, 11, 10, 10, -18, 7, 60, -36, -54, -61, -21, -29, -15, -4, -21, 34, 68, 45, 32, 50, 31, 57, 50, 2, -13, -11, -14, -5, -19, 16, -5, -19, 4, 35, 36, -10, -11, 17, -21, -8, 1, 11, 15, 0, 38, 37, 36, 27, 5, 43, 43, 20, -23, -2, 13, -29, -6, -9, -4, -19, 2, 52, 73, -10, 17, -11, -12, -6, -4, 47, 52, 18, 6, 3, -23, -4, -19, 39, 57, 33, -7, 23, -4, -3, -11, -2, 8, -15, -6, 27, 23, 4, 44, 4, -7, 61, 47, 13, 21, 24, 6, 9, -12, 20, -3, 25, 39, 32, 25, 26, -20, -25, 15, 20, -15, -9, 8, -30, 26, 35, 46, 18, 8, -3, -1, 15, 27, 20, 10, 26, 11, 23, 14, 21, 37, 30, 26, 12, 35, -14, 7, -9, -13, 21, -16, -24, 6, 19, 47, 29, 26, 23, 14, 21, 54, 43, 0, 2, 26, 15, 41, 27, 20, 32, 39, 23, 12, -24, 22, 4, -5, -3, -17, 1, 50, 42, 64, 14, 31, 13, 26, 31, 42, 51, 29, 35, 47, 23, 42, 32, 26, -2, 33, 5, -43, -29, -19, 13, 3, 9, -20, 5, 10, 54, 56, 44, -23, 13, 37, 42, 50, 72, 15, 49, 74, 44, 37, 29, 16, 18, -13, 31, 1, -56, -27, -7, -9, 18, 20, -26, 37, 87, 68, 62, 29, 51, 53, 21, 40, 66, 48, 73, 44, 54, 44, 19, 27, -7, 19, 21, 22, 9, 20, -12, -15, 15, 2, -38, 8, 51, 77, 50, 54, 64, 48, 44, 14, 11, 33, 27, 55, 47, 59, 25, -5, -16, 2, 15, -1, 14, 10, -17, -7, 11, -13, -50, -16, 32, 48, 32, 38, 41, 40, -1, 36, 34, 16, 26, 25, 24, 10, 18, -15, -45, 9, 6, 3, -1, 28, -12, 3, -11, 19, -16, -13, 39, 6, -20, 34, 44, 29, 43, 40, 35, 34, 27, -4, 5, -6, 24, -1, -20, 21, -4, -6, 24, 5, -20, 12, 15, 6, -44, -3, 30, -22, -43, -1, 14, 15, 4, 30, 25, 26, 23, -2, 25, -3, -7, 5, -7, 30, 43, 22, 2, 1, -3, -20, 8, 14, -46, 38, 22, 10, -6, -28, -55, -55, -31, -29, 24, -14, -8, -40, -4, -16, -4, 0, 28, 9, 55, 33, 23, 6, -19, 8, 15, -11, 6, 55, 30, 65, 76, 30, 20, 20, -15, -17, 20, 26, -20, 11, 8, -16, -5, 15, 33, 15, 44, 31, 9, 11),
  32 => (16, 8, -17, -6, 18, 14, -18, 7, 17, 7, -3, 0, 3, -21, 22, 5, 33, 75, 5, -24, -12, -9, 1, 18, 0, 7, -12, 12, -11, 19, 10, -9, -2, -10, 19, 14, -15, 5, -20, -12, -51, -12, 21, 19, 3, -28, 5, 12, 13, 31, 28, -5, -13, -10, -1, 13, -2, 12, -3, 12, 5, -16, 17, 11, 19, -6, -43, -22, 23, 19, 1, -12, 16, 6, -23, -15, 16, 29, 13, -17, 4, -37, 21, -18, 1, 3, 14, 18, 9, 14, -15, 16, -11, -31, 4, 33, -10, -20, -24, 13, 26, -1, 3, 3, -3, -22, -42, -29, 10, 47, -19, -17, 1, 11, 0, 11, -12, 14, 2, -15, -27, -19, -20, -18, -45, -17, -3, 9, -10, -13, -15, 12, 6, -19, -14, 20, 34, 43, 6, -11, -20, 16, 8, -13, -10, 20, -1, -30, -27, 9, 22, -17, -45, 13, 42, 15, -18, -11, 19, -9, -32, 18, -34, 0, -4, 7, -13, 17, -8, -12, 3, 1, -13, -12, -14, 4, -2, 39, 24, -10, -10, 7, 27, 17, -1, -12, -16, 15, 5, -6, -13, -13, -35, -18, -6, -1, 13, -20, 10, 6, 11, -17, -14, 11, -12, -5, -33, -1, 1, 19, 40, 13, -18, -53, -20, -2, 15, 16, 27, 17, -54, 27, -16, -18, -10, -3, 12, -17, 2, 8, -30, 6, -18, -21, -19, -19, 9, 35, 23, 21, -4, -30, -35, 21, 30, 16, 27, 21, -38, -51, -39, -31, 14, -1, 5, 17, 3, -8, 32, 13, 6, 25, 16, -26, 5, 22, 7, 13, 21, -51, -28, -10, 15, -8, 29, 7, 0, -1, -27, -30, 4, 12, -8, -13, -19, 29, 47, 16, 11, 13, -39, -61, -10, -10, 35, 16, 8, -45, -46, 3, 6, 28, 14, 9, 10, 14, 12, 20, 18, -4, -4, -13, -5, -24, 54, 22, 30, 25, -45, -20, 8, 27, 24, 11, -10, -72, -68, -17, 23, -5, 17, 47, 8, 34, 3, 24, -14, -20, -1, -2, -39, -39, 5, 30, 42, -31, -66, -38, 29, 17, 29, 40, -8, -76, -79, -7, 53, 32, 23, 11, -13, 3, 35, 41, 14, -15, -16, -8, -23, -13, 27, 4, 0, -30, -42, -31, 29, 17, 25, 43, -4, -70, -70, -4, 48, 11, 12, 27, -2, 17, 0, 58, -8, 16, 9, -4, -32, 5, 19, 40, -44, -79, -66, -28, 42, 26, 19, 51, -10, -115, -86, -49, 56, 30, 23, 3, -13, -29, 1, 33, -1, 0, -12, -17, 35, 17, 46, 30, -51, -77, -61, 4, 20, 44, -16, 44, -23, -66, -91, -25, 40, 25, -12, 17, -9, -20, -12, 37, -18, -7, 19, 14, 30, 26, 70, 30, -36, -49, -52, -41, 41, 23, 31, 33, -47, -66, -47, -44, 20, 56, 10, 30, 18, 14, -13, 48, -10, 9, 20, -2, -8, -7, 39, 17, -50, -44, -45, 15, 13, 30, 20, 8, -1, -40, -39, -60, 24, 75, 7, 19, 23, 2, 4, 33, -17, 13, 4, 19, -1, 17, 15, -30, -64, -72, -69, 2, 61, 27, 28, 8, -44, -51, -60, -73, 13, 53, 5, 21, 37, 24, -7, 34, 2, 3, -11, -11, -33, -16, 6, -21, -85, -78, -50, 25, 37, 35, 21, 38, -34, -80, -75, -55, 15, 72, 13, 30, 17, 0, -12, 39, 1, 2, 18, 2, -24, -14, -12, -26, -28, -60, -74, 43, 67, 21, 35, 19, -24, -64, -56, -38, 24, 72, 69, 51, 31, -27, 22, 43, 21, 11, 1, -17, -29, -16, -9, -16, -43, -60, -36, 8, 18, 9, -4, 26, -28, -53, -59, -52, -16, 50, 14, 40, 32, -1, 8, 7, 12, 0, 18, 5, -34, -15, 9, -29, -29, -45, -36, 2, 34, 1, 17, -15, -29, -35, -56, -37, 6, 37, 52, 18, 8, -23, 20, -25, -17, 14, -12, -11, -6, -20, 7, -21, -35, -53, -16, 45, 12, 11, 3, 10, -63, -31, -63, -55, -1, 47, 51, 18, 6, -9, 27, -6, -2, 19, 9, 17, -32, -52, -38, -42, -32, -54, 35, 47, 38, 0, 34, -11, -43, -30, -33, -9, -4, 0, 25, 4, 8, -15, -3, -9, 5, -9, 18, -3, 1, -40, -15, -37, -9, -6, 13, 32, 33, 36, -7, -43, -63, -56, -30, -14, -24, -24, 24, 24, 12, 0, -20, -30, 15, 9, -10, 3, 8, -27, -21, -33, -33, -36, 32, 18, 10, 52, 10, -11, -35, -27, -10, -20, 17, -3, 27, -9, 1, 0, -32, -21, 8, -20, 5, 6, -9, 18, -5, -15, 12, 15, 7, -14, 17, 2, -22, 10, 14, -8, -21, -30, -9, -15, -9, 14, -26, -16, -31, -28),
  33 => (-3, 12, 13, -7, 11, -13, 6, 14, -14, 19, 6, 7, -17, -17, -29, -27, -18, -11, 0, -9, -12, 3, -5, 1, 1, -18, -2, -13, 0, -6, -1, -18, -16, -9, 19, -10, -5, -4, 8, 9, 10, -8, -2, 20, 13, 11, 5, 16, -11, -11, -28, 19, 13, -3, -1, 7, 19, 2, 9, 0, -21, 20, -16, -16, -3, -14, 19, -47, -37, 27, 35, 13, 30, 35, 32, 52, 38, 2, 2, -3, 3, 0, -19, 5, -3, 17, 19, 4, 15, -7, 20, 2, 1, -38, -4, 21, 29, 19, -9, -1, -2, -69, 1, 26, -19, 1, -3, -23, -32, -14, -6, -5, 15, 0, 5, -18, -3, -19, 9, -18, -29, -40, 3, -33, -37, -7, -36, -30, -34, -1, 3, -8, -32, -5, -3, -50, -51, 3, 0, 18, -20, -11, -5, 8, 18, 9, 14, -32, -21, -18, -41, -50, -21, 6, -10, 37, 16, 30, 2, 5, -44, -40, -39, -51, -42, -23, -18, 20, -4, 18, 15, -10, 1, -10, -27, -38, -34, -26, -16, 20, 15, -19, 11, 14, 24, 55, 19, -6, -19, -47, -45, -20, -11, -7, 10, -1, 2, 10, -16, 0, -4, 1, -20, -37, -35, -34, 8, 11, 2, 0, 9, 4, 9, 35, 21, -5, -13, 16, -59, -28, 2, -24, 4, 19, 9, -19, -18, 7, 15, -7, -1, -1, -11, 19, 27, 35, -1, 12, 0, -9, 15, 15, 3, 2, 8, -27, -30, -30, 5, -2, 11, -8, 1, -5, 5, -14, 13, 3, 9, 16, 33, 59, 28, 24, 61, 39, 10, -21, 22, 47, 43, 41, 15, 5, -38, -32, -31, 42, 14, 8, 14, 10, -11, 4, 10, -19, -30, 38, 52, 46, 36, 31, 40, 20, -13, -39, 0, 22, 31, -1, 24, 21, -6, -22, 20, 51, -20, -2, 12, -12, -14, 1, -12, -18, -5, 75, 26, 22, -1, 18, 19, 22, -61, -49, -9, 3, 24, -3, 18, 34, 1, -13, 30, 48, -17, -18, 2, -9, 14, -17, -23, 21, -9, 26, 1, -11, -29, -24, -7, -52, -75, -82, -54, -47, -13, -40, -19, -15, -27, -46, 10, 41, -9, -2, 17, 6, 13, -12, 16, -23, -53, -45, -37, -19, -21, -36, -53, -73, -49, -56, -58, -58, -49, -54, -48, -22, -24, -42, -20, 11, -46, -31, -14, 16, -8, -6, -22, -5, -46, -80, -84, -43, -73, -54, -63, -57, -52, -46, -58, -62, -48, -80, -33, -37, -20, -21, -6, 0, -14, -11, -16, 12, -5, -12, -13, -13, -1, -61, -40, -32, -20, 12, 7, 14, 16, -14, 10, -32, -17, -37, -11, -18, -36, -3, -41, -23, 4, -2, -20, -18, -3, 3, 9, 17, -13, -23, -7, 27, 42, 21, 40, 27, 45, 63, 41, 38, 13, 17, -9, 12, 8, 4, -1, -7, 50, -5, 1, -2, -20, -15, 22, -14, -18, -4, 42, 16, 23, 8, -2, 39, 42, 68, 59, 14, 19, 45, 26, 41, 49, 24, 66, 43, 49, 14, 9, -10, 17, -13, 38, 25, -15, 9, 32, 14, -5, 55, 35, 10, 24, 43, 35, 7, 24, 37, 21, 54, 38, 19, 51, 32, 45, 27, 11, -19, -8, -11, 16, 17, 2, 23, 15, 28, -12, 40, 43, 29, 28, 30, 27, 34, 29, 23, 14, 33, 29, -20, 22, 13, 28, 0, 15, -1, 13, 14, 57, 46, 28, 28, 8, 10, 1, 20, 33, 30, 32, 21, 35, 31, 33, 51, -6, -27, 6, -5, 23, 4, 21, 1, 16, 1, 17, -14, 55, 54, -9, 40, -16, -3, -3, -5, -1, 38, -12, 7, 39, 22, 18, 38, 31, -1, 5, 6, 24, 12, 13, 4, -3, -5, -15, -10, 37, 16, -27, -26, -60, -28, -64, 4, 25, 6, -17, -16, 29, 23, 8, 44, 6, 13, 17, 18, 17, 45, -18, 1, -5, 2, 2, 12, 19, -26, -25, -57, -39, -31, -49, 2, 1, -35, -15, -25, 11, -8, 24, -24, -8, -37, 12, 34, 48, 19, 6, 21, 15, 10, 18, -5, -16, -21, -46, -53, -53, -47, -53, -12, -44, -53, -60, -42, -48, -46, -16, -2, -8, -7, -41, -12, 12, 22, 13, 29, -2, 3, 14, 15, 1, 3, -5, -13, -50, -37, -59, 1, 3, 0, -74, -48, -74, -60, -35, 31, -24, -18, -21, -15, -49, -20, -15, 7, 8, 13, 17, -5, -16, 33, 10, -26, -42, -21, -15, -18, 1, -32, -44, -40, -63, -24, -25, -3, -11, -36, -19, -40, -70, -57, -37, 27, -2, 14, 18, 8, -16, 26, 25, 25, 44, 16, 39, -3, -7, -48, -26, -33, -39, -54, -39, 4, -3, 5, -16, -21, -20, -45, -47, 16),
  34 => (-5, 4, -16, 20, -13, -1, -10, -10, -14, -17, -12, 14, -9, 12, 16, 58, -7, -20, 17, 20, 28, 5, 14, -9, 15, -14, 4, -7, -16, -6, 3, 11, -20, -2, -12, 7, -11, -3, -17, 31, 49, 33, 24, 15, -11, -5, 8, 29, 19, 11, 16, -11, -17, -20, -1, 18, 9, -10, 9, 20, -14, 11, 4, -8, 11, 15, 42, 24, 24, 28, 9, -54, -43, -14, 38, 33, 71, 32, -14, -20, 9, 25, -16, -13, 5, 18, -8, 10, 10, 14, 17, 19, -24, 37, 4, 29, 45, 13, -3, -7, 1, 0, 16, 13, 11, 2, -27, -15, 43, 30, 10, -6, 0, -3, -18, 9, 9, -20, -5, -22, 0, 13, 31, 56, 8, -20, -7, 27, -2, 7, -15, 25, 4, -8, -38, -23, 22, 58, -13, -19, -15, 10, -5, -7, 13, -1, -14, 1, -30, -23, -7, 28, -11, -37, -15, -8, 19, -2, -2, 23, 26, -15, -21, -58, 5, 46, 2, -14, -19, -17, 5, 19, -6, -19, -3, 23, -20, -47, 18, 22, -37, -14, -4, 6, 64, 18, -1, 6, 8, 2, -28, -30, 15, 50, 26, 18, -4, 10, -20, 14, 0, 7, 37, -26, -9, 3, 21, 14, -4, -18, -12, 21, 31, 3, 19, 10, 18, 4, -1, -26, 12, 71, 16, -27, 7, -4, -11, -10, -20, 10, 32, -24, 5, 35, 14, -23, -34, -16, -9, 6, 17, 2, -2, 8, 8, -36, -16, -11, 1, 50, 21, -66, 2, -9, -17, 11, 7, -20, 14, -32, 24, 27, 12, -14, -17, -4, -4, 12, 37, 11, 32, 8, -8, 15, 16, 28, 8, 26, 8, -28, -5, 3, -20, 0, 2, -39, 20, 6, 34, 7, 13, -35, -24, 16, 19, 11, 38, 32, -13, -11, -19, -31, 32, -14, -32, 13, 16, 15, 10, 16, -6, 9, -10, -29, -24, -8, 23, 29, 1, -52, -43, -13, 14, -4, 43, 11, -33, -36, -58, -47, 29, -6, -31, -20, 20, 50, -12, -5, 18, -8, 21, 0, -38, 19, 44, 49, -24, -94, -51, 35, 6, 29, -6, -20, -20, -27, -59, -38, 12, 12, -46, -16, 34, 56, -12, -12, -13, -16, -9, -35, -27, -13, 51, 22, -31, -94, -31, 30, 25, 22, 15, -4, -31, -14, -37, -40, -6, 22, -33, -27, 34, 80, -9, -14, -3, -2, -1, -11, 10, 26, 48, -19, -72, -83, -7, 18, 21, 22, 4, -8, -65, -37, -32, -35, 2, 41, 18, -8, 47, 88, 17, -17, -7, -4, -16, -34, 46, 43, 42, -18, -97, -87, 4, 26, 30, 15, -1, 10, -71, -32, -22, -23, 15, 15, -4, -11, -13, 28, -13, 11, 5, -2, -7, -44, 37, 45, 28, -50, -110, -79, 12, 36, 30, 21, 21, 8, -49, -39, 3, -3, 1, 28, 7, -3, -2, -3, 13, -2, 10, -16, 10, 7, 27, 32, -10, -37, -78, -81, 46, 70, 48, -3, 1, -36, -37, -5, 30, 8, -19, 20, 26, 16, 13, -3, -14, -6, -12, 14, -8, -2, -8, 31, -7, -59, -123, -71, 44, 67, 60, 30, 38, -42, -8, -15, 24, 37, -9, 11, 20, -10, -5, -10, -5, 14, 14, -19, -17, -2, 6, 24, -46, -83, -143, -73, 45, 63, 46, 33, 26, -2, -18, -33, 0, -16, -16, -11, 1, -2, -14, -7, 14, 14, 0, -1, 28, 5, 21, 10, -44, -120, -151, -58, 29, 42, 67, 38, -3, -8, -52, -14, 5, 17, -31, 7, 5, -23, 0, -25, 12, 17, 1, 10, 0, 19, 27, 3, -67, -93, -105, -55, 47, 35, 52, 30, 4, -43, -47, -16, -14, 19, -9, 1, 21, 0, 41, -19, -15, -8, -9, 19, -18, 15, 65, 8, -66, -127, -101, -37, 61, 67, 32, 52, 28, 25, 0, -43, -1, -9, -4, 8, -19, 1, 33, 6, 14, -11, 12, -19, -8, -4, 45, 17, -29, -74, -88, -16, 43, 38, 0, 44, 3, -26, -16, -26, -29, -2, -17, -6, -19, 1, -8, 20, 14, 4, -20, 12, -14, -17, -4, -9, -46, -72, -26, 5, -13, 33, 11, 3, 25, 14, -26, -18, 3, -10, 7, 5, -50, -58, -53, 30, 7, -2, 14, -19, 30, 20, -15, -19, -22, -58, -43, -24, 15, 21, 34, -5, 6, 8, 7, -30, -18, -37, -19, 0, -47, -11, 4, 12, 6, -13, 7, 20, 12, 8, -12, -14, -23, -33, -4, 26, 11, -7, 29, -6, 14, 10, -17, -25, -25, -5, -21, -44, 8, 8, 16, -13, -2, 7, -14, -19, 13, 3, 22, -6, 2, -1, -15, 19, 16, -7, -6, -9, -22, -16, -20, -12, -66, -5, -37, -44, 3, -6, 5, 0),
  35 => (10, -17, -1, 17, 10, 9, 12, 15, -6, -13, -14, 15, -11, 6, 16, -10, -18, -40, -12, -44, -12, -19, -2, -16, 1, -10, -8, -19, -18, 8, -10, 4, -10, -14, 20, 5, -11, 6, -5, -14, 0, 35, 0, 14, -7, 3, 6, -12, 5, 3, 21, 21, 3, -6, -6, -3, -17, -10, -6, 16, -3, -3, -20, -8, -4, -17, 19, 1, -9, -11, 1, 19, -7, -9, -22, -15, -1, -16, 22, 34, 15, 20, -18, -15, 7, -5, -12, -6, 13, 5, -2, 19, -14, -54, -29, 7, 2, 13, -6, -12, -7, -36, -50, -21, -21, -16, 17, 39, -11, -18, 20, -1, 9, -14, 3, 14, -8, -12, -20, -12, -41, -20, -11, 31, 37, 38, 18, -10, -33, -31, -38, -23, -37, -41, 5, -8, 2, 35, 19, -14, 8, -3, -8, -13, 11, -4, 8, -40, -8, 47, 37, 36, 25, 33, 14, 33, -1, -14, -35, -33, -23, -36, -17, -6, -12, -7, -8, -9, 2, -7, -15, -18, 2, 16, -33, 2, 6, 12, 38, 15, -30, -33, -11, -22, -53, -19, -44, -39, -51, -20, -22, -16, -7, -13, -10, 20, -6, -5, 5, -2, -19, -2, 22, 2, -10, -11, -20, 16, -32, -37, -36, -40, -27, -14, -7, -1, -30, -8, -23, -22, -16, -4, -10, -10, -14, 3, 19, -14, -19, 17, 21, 18, -35, -77, -39, -37, -39, -32, -13, 23, 2, 17, 4, 7, -13, 13, -16, -30, 15, -27, 3, -2, 17, 15, 5, 7, -10, 7, -33, -39, -73, -51, -25, -11, -2, 2, -12, 26, -13, -21, 21, 37, -27, -19, 16, 8, -3, -28, -4, -8, 10, -9, -19, -14, 14, -8, -35, -28, -67, -50, -32, -19, 13, 7, 14, 17, 9, -52, -50, 2, 25, -29, -17, 28, 1, -8, -12, -10, 16, -9, 11, 7, 17, -23, -14, -24, -2, 3, -32, -43, 18, -29, 9, -9, -45, -34, -19, 29, 6, -11, -19, 24, 25, 14, -15, -17, -4, -13, 20, 6, -18, 11, 31, 28, 17, 8, 10, 9, 12, -13, -16, -61, -44, -61, -34, 7, 20, -11, -9, 12, 20, 7, -16, -13, 9, -10, 2, -19, 23, 26, 41, 61, 41, 22, 6, -18, -34, -50, -41, -74, -78, -71, -41, -8, -9, -9, -36, -8, -10, 8, -27, -27, 5, 18, -12, -2, 15, 31, 20, -13, -2, -16, -12, -46, -46, -75, -45, -59, -82, -48, -53, -47, -4, -42, -33, 13, -4, -7, -25, 5, -15, -14, -13, -16, 3, -1, -44, -54, -4, -14, -53, -76, -34, -66, -19, -32, -51, -24, -11, -4, 1, 0, -39, -18, -28, 3, -45, -9, -13, -11, -6, 17, -15, -8, -52, -51, -25, -29, -50, -55, -58, -52, -58, -80, -23, -1, 14, 2, 22, -35, -6, -7, 4, 10, -10, -3, -17, -2, 5, -3, -6, -11, -47, -39, -17, -35, -49, -32, -52, -65, -33, -30, 31, 12, 20, 23, -7, -9, 4, -4, 8, 30, 25, 16, 10, -9, -20, 11, 38, 44, -55, -55, -29, -40, -64, -17, -13, -30, -26, 6, 58, 44, 28, 7, 1, -18, -18, -12, -20, -16, 43, 15, 17, -17, -18, -12, -19, -20, -34, -41, -21, -30, -35, -2, -2, -16, 14, 26, 49, 29, 31, 30, 31, 20, 21, 10, -24, 13, 42, 34, -15, -15, -8, -13, -20, -22, -51, -7, -26, -45, -51, -24, -29, -3, 10, 41, 27, -8, 17, 55, 43, 30, 49, 28, 19, 35, 33, 39, -10, -16, 10, -21, 16, -17, -7, 0, -8, -28, -38, -16, -18, -7, 9, -6, -30, -16, 4, 21, 39, 11, 22, -13, 17, 26, 28, 60, 8, 1, 1, -14, -5, 8, -13, -13, -3, -22, -23, 10, -27, -22, -10, 14, 10, -25, -12, -34, -2, -4, 20, 12, 21, 35, 8, 32, -2, 11, 13, 15, -3, 25, -25, -13, 18, 2, -8, -7, -23, -13, -10, -12, -5, -28, -35, -18, 12, -7, -33, -11, 5, 35, 12, 13, -6, -20, -10, 19, 14, -8, -5, 7, 8, 16, 6, -26, -25, 4, 12, 10, -3, -50, -6, -39, 20, 10, -20, -26, 6, 13, 6, 51, -16, 0, 18, -1, 14, -1, 0, 15, -11, 11, -4, 5, -36, -19, -21, 19, -34, -45, -54, -15, 1, -1, 2, 3, -26, 1, 14, 23, 7, 2, -10, 20, 19, 12, -10, 10, 3, 1, -21, -4, -5, -25, -34, -8, 2, -35, -28, 7, 27, 7, -14, -14, -30, 6, 39, 48, 20, -9, 15, 20, 6, 20, 18, -3, -22, -16, -12, 6, -5, 0, 21, 33, -6, 4, 8, -2, 25, 23, -29, 4, -29, -39, 23, -3),
  36 => (-18, 14, 13, -6, 1, 11, -2, -9, 17, 0, 11, -20, 16, -16, -10, -31, -31, -39, -56, -50, -30, 8, -12, 17, -15, -13, 18, 17, -12, -5, -8, 9, -14, 14, -14, 5, -1, 17, 15, 21, 62, 21, 47, 10, 44, 30, 33, 32, 27, 33, 57, 27, 18, 9, 6, 2, 3, -1, -20, -18, -15, 20, -21, -14, -9, 34, 4, 77, 57, 36, 59, 46, -31, -17, -29, 0, 14, 19, 16, 11, -11, -10, -8, 18, 17, -6, 3, 19, 9, -8, -17, 16, 46, 3, 15, 21, 69, 80, 33, 2, -13, -46, -37, -21, -23, 1, -17, -13, 4, 37, -20, 1, -12, 1, 19, -10, 9, 12, 6, 18, 5, -43, -22, 28, -3, 35, 22, 2, 14, -20, 14, -8, 10, -15, -12, 9, 9, -10, 2, -19, -13, -8, -7, 8, 4, 9, 47, 4, 26, -22, -32, 18, -32, -3, -1, 12, -3, 15, 24, 6, -19, -9, -22, -19, 26, 28, 13, 7, -10, -14, 7, 11, 5, -17, -9, 66, 71, 10, 24, 34, 20, 55, 18, -18, 7, -1, 12, 19, -24, -22, 4, 11, 24, -10, 12, -16, -3, -4, -6, -14, 5, -16, 65, 98, 51, 34, 59, 31, 59, 32, 14, -2, 26, 11, 6, 8, 5, 6, 16, 2, 7, 11, -2, -35, -12, -7, -17, -19, 9, -4, 70, 68, 44, 25, 80, 55, 40, 36, 24, 47, 4, 29, -3, -5, 26, 13, 3, -18, 33, 27, -10, -25, 10, 21, -17, -3, 13, -9, 58, 42, 31, 34, 55, 30, 9, 27, 34, 31, -7, 24, 27, 22, 8, 39, 17, 31, 1, 22, -14, -22, -7, 12, -13, -11, 19, 12, 13, 24, 27, 26, -4, 3, -8, -17, 11, 13, 27, -1, -25, -43, -2, 20, 34, 27, 20, 6, 3, -10, -3, 14, -18, -2, -15, -52, 31, -14, 2, 37, -9, -21, 0, -13, -7, 2, -4, 1, -47, -16, -13, 18, 21, -9, -13, 24, 17, -53, 8, -10, 5, -14, -27, -61, 31, -3, 29, 24, 20, 12, 35, 27, 15, 7, 11, 15, -14, 32, 22, 37, 45, 31, 24, 38, 37, -19, -8, 18, 16, 17, -3, -30, 48, 23, 45, 37, 43, 48, 29, 14, 39, -6, 23, 29, 25, 68, 91, 75, 61, 31, 42, 48, 41, -12, 16, -6, -11, 4, -4, -5, 27, 45, 50, 46, 43, 29, 44, 14, 44, 57, 63, 63, 65, 58, 90, 104, 62, 40, 60, 66, 53, 8, -14, -3, 15, -15, -18, 13, 13, 31, 26, 56, 67, 42, 64, 20, 34, 71, 79, 54, 69, 88, 89, 62, 78, 67, 55, 39, 37, 9, -3, 1, 20, 5, -17, 14, 39, 34, 18, 8, 78, 84, 39, 37, 39, 50, 49, 59, 85, 60, 33, 60, 68, 34, 23, 1, -29, 37, -3, 5, 4, -6, 31, 10, 43, 24, 42, 34, 51, 37, 50, 44, 61, 38, 44, 68, 86, 38, 46, 28, 36, -4, -3, 26, 5, 23, -20, 20, 20, 20, 22, -27, 9, 2, 39, 18, 37, 51, 52, 57, 32, 15, -21, -1, 48, 45, 26, 38, 51, 10, -10, -17, 38, 55, -9, 13, -17, -11, 25, -25, -15, -11, 14, 56, 28, 39, 28, 33, -5, -32, -13, -5, 29, 39, 35, 67, 59, -3, -12, -24, -6, 1, -15, 18, -18, 0, 7, -15, 7, -13, 12, 10, 63, 30, 6, 24, 30, -25, -5, -7, -9, -5, 25, 25, 58, -4, -24, 12, -8, -39, 20, 10, -12, 17, -9, -28, 3, -32, -29, -15, 6, 15, -5, -22, 21, 8, 33, 18, 17, 49, 14, 25, 16, -13, 9, 8, -4, -23, -20, 6, -16, 0, -39, 15, 21, 18, 8, 5, -4, 5, -8, 12, -3, 7, -25, -5, 7, 17, 20, 17, 22, -33, 2, -5, -13, -50, -17, -20, 18, 12, -39, -21, 9, 40, -4, 4, 13, 40, 12, 39, 17, 25, 47, 18, -1, 14, 44, 29, 15, -20, -9, -14, -25, -43, -3, 14, -10, 20, -15, -37, -20, 16, -7, 10, 62, 34, 8, -7, 21, 41, 35, 1, -23, 5, 11, 15, -14, -40, -5, 22, 3, -27, -11, -4, 16, -2, -54, -34, -7, 13, 26, 34, 57, 12, 3, -24, 32, 48, 25, 43, 22, 14, -7, -13, -45, -38, -12, -5, -24, -49, 15, 17, -19, -5, -6, 15, -22, -28, -11, 7, 47, -10, 21, -14, -14, 15, 14, 13, 23, 36, 53, 41, -13, -34, 11, -27, -49, -48, -3, 10, 15, 15, -20, 38, 19, 59, 63, 41, 35, 29, 37, 26, 50, 52, 31, 44, 24, 9, 48, 18, -30, -9, -5, -14, -44, -52),
  37 => (-3, 0, 8, 9, -3, -9, 8, 10, -16, -14, 9, 20, -4, -8, -3, -7, 17, -10, 16, 23, 17, 16, -9, 12, -12, 16, -2, 13, -19, -19, -14, -6, -20, -10, 18, -6, -18, -12, 0, 17, 5, -16, -45, -29, -2, 12, -24, 2, -8, -10, -14, 4, -4, 14, 5, -9, 5, -1, 11, -20, 2, -18, 20, 15, 6, -12, -20, -34, -25, -66, -59, -25, -12, -31, -63, -26, -14, -4, -22, -27, -14, 15, 5, -13, -16, -3, 9, -15, -8, 9, -15, -2, 5, -24, -45, -65, -50, 13, 7, 14, -17, -8, 0, -35, -10, -16, 25, 2, -12, 27, 18, -14, -5, 8, -7, 12, 14, 15, 8, -20, -8, -68, -79, -75, -30, -5, -17, -19, -24, -26, -39, -39, 7, 14, 27, 34, 48, 15, -13, -19, 14, 13, 1, 16, 17, 12, -17, -28, -63, -95, -75, -70, -39, -26, -43, -4, 2, -13, -65, -39, -38, -1, 21, 18, 30, 46, 14, 2, -2, 19, -14, -19, -2, -9, -21, -39, -110, -106, -86, -50, -41, -25, -32, -24, -8, -1, -2, -38, -40, -28, 23, 19, 24, 67, 17, 8, -4, 2, -11, 6, -2, 20, 15, -33, -67, -46, -35, -24, -10, -15, 25, -1, 23, 19, 5, -20, -52, -56, 3, 14, 19, 54, 3, 4, 4, 17, 2, 19, 18, -13, 11, -16, -18, 0, -23, -17, -11, -34, -1, 2, 12, 26, -14, -41, -36, -57, -37, 11, 30, 37, 20, -18, 3, 10, 11, 11, -19, 18, 24, -27, -16, 21, -10, -35, -45, 11, 47, 21, -11, 7, -30, -2, 2, -49, -27, 4, -18, 37, 37, -21, -8, 1, 15, -4, -18, 3, 32, 2, 31, 46, -14, -16, -29, -22, 26, 17, -24, -19, -21, 11, -10, -23, -7, 6, -10, -8, -1, -4, -7, 6, 13, 16, -15, 58, 69, 13, 53, 44, 39, -6, -33, 13, -8, 19, 2, -20, 5, -6, -3, -19, 0, 1, -18, -31, 8, 28, -15, -12, -17, 1, 17, 54, 65, 57, 74, 48, 14, -28, 33, 12, 24, 21, -23, -9, 41, 18, -11, -18, -13, -21, 4, 1, 3, 55, -19, -8, -11, -16, -10, 48, 14, 32, 34, 22, 40, 27, 67, 44, 59, 43, 46, 28, 48, 29, -11, 6, 9, -13, 43, 4, 15, 56, -8, 3, 5, 0, 42, 34, 22, 44, 37, 56, 77, 48, 67, 66, 50, 60, 56, 27, 36, 33, 9, 4, -14, 20, 33, 0, 35, 33, 17, 5, 9, -19, 31, 25, 42, 39, 14, 1, 25, 50, 29, 48, 54, 57, 46, 37, 36, 11, 14, 26, 11, 17, -1, 12, 6, 42, 12, -9, 19, -4, -19, 52, 25, 9, -2, 17, 8, 2, 19, 8, 17, 36, 63, 53, 24, 4, 17, -2, 37, 27, 6, -3, 23, 63, 4, 19, 1, 3, 51, 23, 7, 13, -24, -1, 0, -6, -9, 30, 34, 38, 34, -18, 27, -3, -7, 7, 2, 28, -19, -26, 12, 74, -9, 17, 13, -18, 33, 44, -23, 8, -24, -39, -46, -89, -43, -11, -6, -15, -14, -20, -25, -20, -9, -15, 12, 19, -2, -9, 16, 92, 15, -4, 8, -20, 16, 9, -33, -45, -71, -106, -146, -99, -45, -47, -13, -19, -34, -42, -42, -27, -39, -8, -26, -16, -29, -44, 21, 53, -9, -5, 11, 17, -30, -62, -69, -69, -76, -96, -140, -58, -34, -2, 2, -17, -48, -43, -35, -45, -36, -51, -47, -23, -22, -40, -18, 45, -1, -16, -5, -1, -23, -66, -61, -73, -88, -132, -129, -74, -10, -5, -28, -4, -43, -59, -32, -35, -28, -35, -25, -13, -2, -79, -21, -8, -15, 3, 6, -17, -20, -43, -54, -49, -62, -101, -80, -54, -4, -24, -7, 35, -28, -20, -19, -13, -43, -21, -23, -19, -10, -33, -22, -3, 18, -21, 17, -20, -1, -51, -61, -48, -55, -54, -99, -51, -14, -44, -1, -4, -42, -43, -18, -31, -45, -34, -34, -11, 0, -1, -5, 17, 7, 15, 12, 17, 19, -22, -40, -37, -1, -18, -55, -29, 26, 10, -13, 2, -37, -17, 7, -27, -45, -11, -59, -25, 22, 12, -10, 12, 0, 1, -18, 4, 28, -5, -26, 1, -12, -17, -15, 15, 29, 33, 6, -4, -11, 32, -5, -6, -20, -52, -16, -15, 30, -2, -9, 11, 0, 18, 14, 14, -2, 20, 50, 8, 2, -8, -38, -2, 6, 25, -35, -27, -34, 1, 17, -33, -41, -25, 3, -16, 37, 20, 22, 13, 17, 10, -20, -5, 12, 14, 5, -19, 10, -19, -2, -8, -12, 24, 43, -21, -42, -31, 44, 43, 15, 32, 36, 28, 37, 88, 56, 56),
  38 => (19, -19, -4, -5, -20, 7, -14, -18, -12, 20, 13, 13, -17, 7, -8, -23, -50, 29, 13, 32, 14, 7, -22, 8, 0, -1, -18, 16, -13, 8, 14, -12, -6, 3, -3, 17, 7, -12, 13, 2, -48, -1, -12, -29, -37, -16, -45, -23, 17, 33, -17, 10, -11, 8, -3, 19, -2, 21, -8, 2, -1, -5, -9, 6, 7, 8, -9, -41, 8, -1, 18, -1, 15, 20, -16, 22, 47, 3, -19, 15, -4, -8, -3, 20, 11, 8, 4, 15, 4, 5, 12, -7, 14, -24, 1, 44, 73, 49, 30, 52, 6, -5, -18, 33, 21, 11, -30, -43, -27, -22, 4, -13, -3, -11, -14, -7, 2, -16, 15, -15, -9, -3, -7, 18, 43, 41, 41, 32, 28, 57, 58, 24, 27, 28, 8, -18, -34, 15, 8, -5, 9, -19, 3, -17, 10, -15, 10, 12, -28, -39, -54, -17, -1, 68, 41, 11, 62, 64, 44, -7, 42, 17, 63, 46, 14, -34, -11, -11, 0, -19, 9, -17, 6, 11, 14, -28, -43, -29, -20, -19, 5, 40, 13, 17, 46, 37, 7, 24, 18, 42, 48, 77, 50, -7, 15, 11, 3, -9, 4, 6, 14, 19, -36, -31, -67, -43, -45, -52, 1, 12, 24, 22, 39, 43, 44, 33, 37, 65, 39, 71, 51, 30, -8, -30, -13, 7, 17, 9, -10, 11, -43, -51, -44, -58, -70, -67, -53, -26, -71, -67, -10, 42, 55, 23, 24, 14, 7, 51, 58, 65, 0, 4, -5, 17, -20, -11, -11, 3, 12, -57, -7, -35, -24, 21, 4, -38, -70, -74, -38, 25, 56, 32, -6, 23, 24, 47, -2, -17, -23, -59, 6, 17, -6, -3, -19, -15, -53, -32, -26, -16, 25, 21, -40, -73, -43, -23, -19, 15, 37, 36, 4, -4, -11, 34, -12, -20, -21, -62, 11, 17, -14, -7, -1, -11, -68, -33, -14, -47, -42, -70, -66, -102, -31, 2, 21, 49, 1, 24, 27, -19, -11, 7, 4, -45, -23, -40, -17, 3, 12, -1, -13, 13, 1, 39, -27, -33, -28, -11, -41, -9, 22, 28, 38, 16, 4, 4, 13, -33, -6, -10, -20, -48, -30, -66, -9, -18, -11, 19, -14, -2, 25, 7, -72, -62, -32, 19, 10, 36, 25, 76, 31, -38, -51, -4, -5, -30, 15, 16, -16, 11, -30, -51, -10, 10, -2, 14, 15, -28, -17, -45, -73, -45, -9, 7, 24, -8, 5, 25, -19, -22, -51, 15, -19, -40, 25, 13, -18, -7, -29, -3, 18, 2, 9, -1, 57, -14, -6, -20, -44, -29, 13, 18, 30, 18, -4, 6, -28, -18, -37, -4, -2, 15, 29, -8, 35, 11, 6, 20, -14, 13, -7, -12, 27, -1, 50, 34, 51, 8, 71, 38, 24, 1, 15, -15, 0, -1, -20, -17, -20, -12, 10, 4, 26, 39, -29, -26, 2, 12, 12, 13, -9, 40, 60, 70, 52, 42, 41, 30, 41, 26, 43, 11, 21, 3, 2, -22, -34, -25, 31, 8, -1, 26, -22, -40, -15, -8, -15, -2, 26, 86, 69, 47, 8, 34, -8, 35, 7, 32, 25, -5, 5, 12, 34, -12, -45, -36, -30, -15, 24, 38, 6, -59, -10, 11, -9, 7, 42, 34, 74, 60, 7, 43, -9, 15, 29, 32, 15, 11, -26, -7, 14, -13, -79, -89, 0, -16, -8, 54, 2, -34, -12, -17, -1, 7, 43, 32, 69, 37, 41, -3, -1, -30, -26, 32, -8, -1, -28, -39, -8, -20, -54, -30, -1, -10, 5, 27, 1, -20, 19, -10, 21, -15, 6, 5, 33, 28, 24, 16, 5, -18, 11, 12, -24, -8, 43, -4, -30, -32, -29, 17, 11, 1, 3, 21, -40, -6, 10, -16, 12, 18, -39, 5, 36, 39, 41, 70, 70, 16, 51, -25, -50, -7, 8, -22, -31, -35, -32, 29, 65, 37, 1, 18, -36, -3, 11, 5, 13, -11, 4, 10, 16, 48, 15, 49, 23, -21, -27, -70, -88, -44, -47, -23, -15, 1, 34, 26, 32, 16, -8, -16, -3, 1, 18, 12, 5, -18, -11, -3, -12, 20, -20, 2, 7, -33, -26, -78, -73, -37, -3, -32, -21, 17, 33, 37, 23, -6, -19, 6, 6, -12, 7, -10, -4, 4, -27, 5, 15, -3, -25, 14, 19, -62, -21, -55, -76, -76, -50, -38, -35, -5, 13, 23, 8, 21, -22, 5, -10, 12, 3, 20, -4, 7, -10, -1, 7, -16, -8, -27, 2, -40, -21, -69, -74, -88, -81, -42, -25, -48, -23, 6, 4, -10, -56, -17, 16, 21, 12, -20, 6, 15, -13, -17, 5, -6, -36, -2, -11, -21, 16, -33, -32, -52, -39, -58, -38, -16, -40, 7, -21, -10, -24, 1, -15, 19),
  39 => (-20, -7, 6, -16, 5, 10, -3, -11, -20, 4, -10, 11, 18, 9, 21, -2, -20, -9, -44, -7, 3, 7, -20, -10, 15, 9, -14, -8, 1, -8, 14, -17, 19, 1, 12, 13, -19, -17, -14, 3, 2, 28, -4, 11, 0, -13, -19, -11, 20, -31, 0, 14, -2, -12, -17, 1, -2, 15, 14, 5, -10, 2, -10, 13, -5, -10, -1, 21, 42, 59, -14, -44, -96, -91, -19, 25, 29, 31, 38, 52, 25, 11, 19, 7, -15, 1, 1, -3, -4, -9, 11, 16, -5, 42, 13, 19, 1, -14, -60, -57, -76, 8, 17, 49, 7, -2, 3, 7, -33, -24, -19, 20, 17, 3, 19, -2, -6, -20, -5, 8, 35, 6, -17, -17, -8, -5, -18, -38, -4, 17, 41, 48, 27, -11, -17, -22, 3, -20, -9, 4, -15, -14, 0, 17, 5, -2, -2, 23, -14, 16, -28, -42, -34, -70, -79, 8, 6, 29, 30, 22, 0, -16, -15, -34, 12, 4, -5, -18, 19, -4, 11, -20, -15, 7, -15, -31, 14, 2, -31, -42, -58, -84, -68, 42, 19, 24, 14, 22, 35, -5, -34, -16, 40, 2, 1, 20, 4, 0, 13, 11, 5, -16, -4, -29, 23, 10, -20, -43, -97, -123, -41, 38, 35, 28, 25, 31, 15, -25, -34, -49, 8, 42, -7, -12, -11, -14, -16, -17, -15, -19, -1, -44, 33, -2, -32, -72, -110, -109, -39, 2, 32, 31, 42, 29, 11, -48, -22, -33, 4, 31, -11, -38, 18, -16, -8, 9, 17, -2, -21, -30, -16, 2, -37, -62, -86, -59, 10, 32, 13, 36, 48, -11, 8, -67, -36, -17, -18, 11, -5, -29, 8, 9, 9, -15, -7, -7, -52, -14, -5, -14, -55, -58, -67, -16, -21, 29, 32, 23, 48, 26, -40, -49, -35, -21, -24, 13, -4, 2, -3, 19, 20, -14, 8, 8, -36, 9, 14, 5, -24, -18, -28, -28, 9, 9, 19, 14, 18, -21, -6, -34, -35, 25, -13, 1, 44, -31, -19, 2, -20, -9, 3, -30, 5, 31, 28, 17, -19, -47, -21, 3, 2, 10, 10, -15, -14, -14, -40, -40, -43, 1, -26, 17, 39, -14, 20, 11, 17, -12, -2, 43, 31, 29, 60, 43, -38, -66, -12, 12, 16, 41, 21, -7, 11, -19, -21, -34, -6, -7, 14, 30, 62, -19, 11, -11, 12, 1, 16, 24, 59, 57, 76, 15, -74, -86, -23, 31, 23, -8, -11, -25, -3, -32, -18, -7, -14, -9, 9, 51, 35, 9, -14, 5, 18, 20, -23, -3, 17, 40, 78, 4, -75, -99, -50, -7, 2, -11, 13, 4, -15, -33, -14, 8, 9, 8, 10, 10, 25, -5, 13, 11, -15, -6, 2, 10, 54, 45, 55, -5, -63, -48, -20, 25, -9, -24, 1, 8, -17, -37, -24, 22, 15, 17, -10, -2, -40, -18, 14, -16, -5, 19, 34, 14, 44, 54, 64, 16, -28, -55, -38, 28, -2, 14, -12, 14, -30, -7, 1, 8, -4, 22, 11, 7, 7, -44, 19, 7, 7, 16, -31, -2, 46, 46, 83, 59, -39, -79, -39, 23, 32, 12, 19, 19, -23, -19, -1, 3, -49, 17, -10, -24, -45, -90, 0, -13, -2, 8, -16, -45, 19, 60, 75, 44, -17, -56, -13, -8, 11, 34, -3, 8, -21, -14, -31, -37, -10, -20, -7, 6, -47, -56, 13, 4, -17, -3, -12, -25, 18, 63, 13, 32, 4, 4, -1, -2, -1, 7, 11, -16, -8, -6, 17, -12, -18, -6, -26, -32, -9, -60, 11, -13, 17, -11, -16, 18, 22, 23, 43, 24, 5, 11, -10, 13, -16, -10, -24, 18, 8, 51, 14, 10, -11, 10, -28, -9, -62, -74, 14, -19, -19, 9, -48, 43, 18, 23, 23, 51, 22, 38, -31, -16, 17, 7, 20, -3, 46, 16, 25, -20, 4, 5, -12, -9, -50, -55, -18, 20, 11, 16, -15, -5, 19, 15, 16, 39, 27, 14, -51, -31, -13, -16, 33, 24, 21, 20, 0, -15, 5, -27, -35, -64, -59, 26, 16, -9, -19, 21, 11, -38, -33, -19, 15, -12, 7, -1, -17, -27, -63, -34, -7, 33, 52, 15, -20, -40, -23, -12, 19, -12, -44, 1, -11, 14, 13, -13, 18, 6, -41, -11, 10, -7, 9, 13, -91, -66, -40, -34, -10, 12, 27, 14, 21, -10, 0, -1, 0, -13, -10, -34, -14, 13, -1, -12, -6, -15, -9, 6, 13, 39, 30, -11, -46, -58, -80, -26, -13, 3, 12, 8, 34, 19, -25, -15, -25, -24, -1, 26, -9, 4, -3, -8, 19, -15, -15, 19, 35, 16, 11, -17, -18, -62, -44, -33, -34, 0, -5, 35, 17, -5, -15, -42, -51, -2, 47, 6),
  40 => (7, 7, 6, -15, 14, -17, -18, 14, -14, -5, -17, -1, 16, -20, -1, -19, -28, -49, -34, -5, 40, 12, -1, -10, -9, -5, 17, -18, 18, -4, -11, -7, -12, -7, 11, -3, -17, -7, 41, -18, -12, 25, 19, -27, 18, 5, -39, -7, 10, 12, 34, -13, -17, -18, 17, 19, 18, -20, -14, 6, -14, 12, -2, 8, -1, 13, 9, 12, 5, 7, 13, 36, 22, 28, -2, 18, -17, 5, -19, -23, -57, -24, 11, 14, 18, -13, -4, 7, 10, 8, 6, -19, 14, 4, -19, 40, 37, 73, 41, 50, 38, 17, 35, -5, 19, 2, 4, 4, -41, -23, 15, 14, -19, -1, -7, -9, -3, -10, -2, 61, 11, 46, 68, 43, 53, 52, 49, 49, 36, 22, -7, -4, -20, 18, -13, 15, -11, -25, 14, -3, 1, 7, 3, -11, -16, 10, 38, 30, 43, 137, 119, 92, 62, 64, 48, 56, 24, 51, 0, -15, -11, -5, 21, 3, 34, 14, -2, 6, -10, -8, 0, -19, -12, 17, 23, 20, 29, 65, 64, 60, 39, 9, 20, -25, 8, 37, 7, 24, -25, 2, -10, 19, 5, -24, -3, 3, 16, -6, 8, -1, 15, -12, 13, 47, 31, 46, 50, 68, 32, 36, -3, 20, 31, 40, 32, 45, 24, 40, 25, 34, 0, -59, -5, -26, -15, 5, -1, -7, -21, 1, 32, 69, 71, 40, 78, 85, 40, 49, 43, 38, 46, 14, 35, 44, 30, 35, 29, 20, -33, -83, -60, -2, -12, -4, -7, -11, 18, -12, 65, 46, 72, 28, 51, 22, -4, -1, 9, 23, -6, -1, 45, 19, 1, 51, 82, 19, -60, -88, -55, -45, 11, 3, -20, 13, 8, -34, 33, -3, -26, -21, -24, -19, -17, -27, 9, -16, 28, 22, 28, 61, 10, 33, 37, 34, -22, -50, 5, -30, 5, 10, -11, -1, -8, -33, -35, -82, -97, -97, -65, -80, -26, -22, -19, -5, 26, 31, 52, 50, 10, 41, 57, 16, -28, -51, -34, -52, -1, 14, 9, 9, 31, -69, -42, -84, -94, -85, -87, -63, -36, -13, -3, -34, 26, 23, 39, 35, 10, 6, 65, -10, -3, -57, -15, -69, -13, 1, -15, 14, 13, -26, -76, -92, -44, -68, -40, -33, -17, 8, 2, 14, 10, -12, -3, 9, -7, -14, -20, -23, -59, -41, -81, -38, 5, -13, 1, 7, -20, -30, -24, -19, 47, 19, 3, -3, 3, 26, -23, -8, -9, -26, -15, -6, -3, -16, 19, -13, -35, -51, -73, -55, -5, -8, -1, -15, -12, 12, 20, 37, 63, 26, 25, -4, 6, 14, 1, 30, 10, -25, 8, 9, -27, -26, -6, -10, -40, -14, -84, -46, -7, 5, 13, -15, -3, 21, 42, 58, 73, 56, 60, 36, -23, 15, 4, 29, 43, 15, 42, 28, -13, -10, -1, -11, -45, -23, -74, -18, -9, -17, -4, 15, -9, 38, 41, 37, 51, 28, 22, 29, 8, 26, 45, 63, 23, 16, 26, 13, 3, -19, 11, -17, -49, -74, -47, -26, 20, -8, 9, -4, -13, -10, -4, -8, -24, -30, -3, 10, -6, -8, 18, 36, 8, 21, 12, 1, -12, -18, 7, 22, 13, -41, -32, -47, -8, 16, -19, 8, -11, -8, 5, 2, -5, 8, -3, 25, 5, -18, 3, 12, 4, -11, -13, 3, -15, -3, 22, 24, 20, -31, -10, -47, -17, -14, -2, 17, -26, 10, -9, -1, -14, -21, 38, 6, -30, 0, 35, 12, -20, 11, -6, -20, -9, 12, 8, -2, -20, -62, -10, -9, 13, 15, 0, 11, -13, 45, 1, -9, 25, 32, 55, 68, 31, 36, 40, 15, 10, 31, 45, 22, -23, -5, 16, 23, 20, -16, -21, -14, -14, 3, 20, -17, 0, 39, 39, 0, 25, 7, 45, 63, 37, 52, 40, 0, 7, 40, 36, 19, -12, -9, -4, 37, 26, 7, 10, -45, -7, -14, 8, 16, 8, 27, 4, -12, 17, -3, 23, 15, 36, 34, -2, 21, 24, 50, 36, -13, -19, 15, 38, 40, 17, -18, 26, -11, 20, -1, 0, 16, -18, 17, 2, -7, -8, 15, 2, 21, 61, 23, 38, 44, 42, 49, 27, 34, 26, 29, 14, 72, 40, -10, 12, -30, -7, -6, -17, -14, 17, -16, 16, -12, -8, 22, 21, 29, 42, 67, 59, 49, 27, 58, 45, 61, 7, 17, 24, 35, -54, -14, -16, -36, 10, -6, 10, 9, 2, 21, -2, 12, -9, 17, -6, 5, 35, 0, 32, 28, 55, 32, 55, 20, 18, 22, 12, 18, -27, -10, -32, -65, 6, -14, 20, 17, 4, -15, -11, 5, -34, 6, 30, 44, 30, 6, 37, 45, 45, 42, 41, 38, 19, -3, -3, -7, 23, -28, -50, -11),
  41 => (2, 6, -7, 9, -16, -4, 0, 10, -12, 20, 2, -5, 19, 11, -3, -19, -40, -52, 16, 34, 11, -15, 15, 12, -1, -18, -1, -12, 13, 0, -5, -9, 3, 10, 10, 4, 20, -2, -16, 13, -14, 1, -31, -25, -28, -18, -15, -13, 3, 5, 13, -16, 0, -16, 5, 6, 8, -18, 9, 17, 11, -18, -17, 17, 6, -17, 13, -9, -56, -36, -15, -38, -14, -1, 12, 2, 4, 8, 31, 25, -5, -11, 17, 12, 3, -5, 17, 8, -11, -19, 3, -15, -3, 6, -16, -26, 26, 46, -9, -5, -2, -17, -10, 1, -17, 4, -5, 68, -9, -4, 8, -5, 5, -8, -10, 17, 19, 8, 16, 10, -13, -2, -26, -6, -16, 7, 11, 2, 10, 0, 35, 26, 15, 2, -10, 27, 21, 28, 15, 18, 14, -11, -6, -19, -18, -20, 9, -3, 12, -20, -15, -50, -27, 8, 31, 17, 42, 41, 47, 40, 25, 31, -3, 11, 50, -29, 18, -12, -12, 20, 7, 6, -15, 5, -6, 13, -24, 19, -26, -45, -39, -11, 14, 16, 48, 46, 17, 33, -3, -7, 15, 22, 50, 21, 1, -15, -1, 12, -4, -1, -18, -5, 7, -17, -30, -28, -42, -71, -88, -49, -39, 3, 38, 33, 42, 44, 37, -7, 24, 35, 60, 12, -7, -12, 11, -8, -13, -13, 17, 0, -12, -31, -10, -67, -57, -26, -63, -90, -26, -23, 56, 73, 58, 32, 46, 16, 25, 38, 2, 15, 2, -6, -9, 14, 0, -1, -11, -7, -13, -59, -55, -29, -39, -46, -76, -65, -14, -28, -20, 24, -6, 42, 9, -10, 17, 33, 0, 18, -10, -9, -14, -4, 0, 18, -18, -10, -1, -35, -33, -19, -38, -51, -48, 3, -25, -17, -11, 24, -3, 21, -11, -37, 13, 28, -11, 2, 0, 22, -15, 4, -17, -19, -8, -19, -14, -33, -35, -19, -46, -28, -12, -42, -50, -13, -9, -6, 20, 7, 8, 9, -2, -5, -20, -27, 14, 12, 15, 1, -15, 4, 4, -7, -20, -51, -56, -29, -36, -50, -54, -71, -55, -18, 2, 12, 8, -1, -26, -25, -15, -33, 0, -30, -12, -40, 1, -13, -4, -10, -5, -11, -29, -48, -57, -80, -98, -91, -85, -79, -20, 18, 8, 12, 18, 7, -14, -14, -16, -35, -14, -10, -24, -8, -3, 12, 1, -15, -20, -23, -68, -90, -102, -93, -122, -107, -74, -25, 29, 59, 38, 31, 3, -12, 0, -21, -29, -3, 0, -11, -52, -21, -18, 8, 9, 10, -11, -18, -59, -106, -92, -89, -38, -31, -3, 10, 56, 73, 36, 17, 6, 14, -17, -10, 9, -52, -50, -35, -27, 6, -20, -15, 7, 7, -17, -23, -36, -91, -42, -13, -9, 9, 9, 17, 71, 47, 63, 7, 1, -3, -3, 23, 22, -16, -30, -20, -34, -7, 14, -11, -1, 19, 12, -13, -83, -48, -5, -20, -8, 28, 25, 59, 52, 64, 48, 18, 11, 28, 10, 4, 14, -10, -8, -11, -25, -14, 18, 18, -9, 8, -4, -68, -66, -2, 1, 9, 39, 16, 16, 33, 80, 73, 46, 8, 20, -11, 17, -2, 10, -15, 1, -20, -27, -28, 19, 20, 14, -2, -22, -85, -33, 1, 2, -25, 3, 6, 18, 24, 56, 61, 62, 19, 32, 22, -14, 18, 1, 6, -4, -11, -20, -4, 4, -6, -19, -15, -2, -52, -10, -1, 3, 12, 8, 7, 4, 16, 44, 25, 23, 28, 18, -4, -10, 2, 11, 20, 12, 16, 25, 18, -7, 9, 18, 7, -18, -8, 8, 4, 30, 27, 63, 67, 35, 41, 17, 22, 2, 12, 23, -3, -5, 2, 14, -2, 20, 25, 47, 20, 20, 4, -2, -2, 12, 30, 42, 14, 40, 37, 36, 43, 26, 8, 11, -5, -46, 5, -13, -11, -37, -2, 2, 21, 5, 13, 6, 43, -10, 18, -11, 2, 4, 71, 53, 52, 39, 34, 33, 23, 29, 32, -1, -43, -20, -38, 12, -46, -38, -13, -41, -12, -8, 19, 13, 44, 9, 13, -2, 0, -14, 73, 37, 19, 11, 33, 20, 14, 38, 15, 13, -31, -2, -18, -41, -44, -57, -36, -18, 1, -22, -43, 14, -24, 14, -20, -6, 2, -27, 17, 30, 23, 21, 49, 33, 31, 4, -4, -9, 13, 8, -18, -39, -32, -48, -54, -35, -19, -47, -24, -36, -51, -9, -10, 20, 5, -7, -16, 14, 2, 12, -6, -6, 0, 31, 2, -9, 22, 0, -10, -23, -24, -40, -4, -13, -37, 16, 2, 15, -9, -13, -3, -14, -9, 9, -25, -37, -34, 4, -26, -16, -30, 28, -2, -16, -17, 2, -31, 10, -25, -21, -41, -71, -21, -8, -8, -13, -7),
  42 => (1, 15, -13, 11, -5, 4, -6, 12, -3, 10, -1, 20, -10, 11, -4, 20, 12, -12, 4, 10, -7, 6, -3, -15, -21, 6, 12, -8, -19, -1, 4, 5, 13, 4, -4, -14, -7, 20, 13, -8, -6, 12, 2, -30, -15, 5, -21, -10, 55, 6, -8, -3, 7, -20, 9, 2, -3, -4, 19, 6, 20, 2, -5, 12, -12, -14, -1, -4, 2, -1, -12, -74, -79, -64, -31, -28, -22, 24, -17, -20, 14, -16, -16, 17, -4, 17, 14, -12, 3, 16, -11, -4, 14, 7, -13, -36, -56, -11, -9, -25, -12, -10, 12, -1, -26, -17, 0, 20, -8, 3, -15, 9, 18, -7, -8, -2, 18, -5, -14, -16, -13, -61, -109, -128, -48, -26, 33, 32, 27, 12, -9, -47, -38, -16, 37, 26, 7, -9, -7, 12, -1, 4, 9, -17, -4, -3, -17, -38, -26, -98, -169, -110, -27, 16, 30, 56, 23, -13, -59, -38, -67, -55, 49, 44, -17, -18, -11, 10, -3, 7, -9, 8, 4, 0, 7, -26, -4, -104, -92, -64, 10, 48, 50, 52, 13, -40, -89, -53, -49, -71, -24, -2, -29, -23, -6, -6, -2, 11, 19, 17, -5, 7, -33, -37, -8, -101, -85, -29, 1, 66, 49, 39, -44, -33, -86, -76, -52, -87, -52, -35, 7, -44, -15, 18, -4, -13, -19, -11, -18, 16, 0, -30, -52, -119, -80, -21, 22, 50, 16, -54, -57, -39, -43, -56, -47, -117, -70, -38, -11, -37, 3, 15, 9, 17, 17, -16, 14, -16, -17, -8, -25, -74, 0, -2, 15, -5, -21, -25, 13, 14, -1, -22, -22, -28, -26, -1, 19, -14, 11, -19, 2, -15, -5, 9, -6, -17, -23, 27, -28, 6, 31, -6, 24, 17, 11, 6, -9, -22, 3, -11, 0, -10, -1, 8, 41, 26, 32, 13, -16, -16, 11, -20, 17, -61, 14, 29, -8, -6, -12, 2, 8, 63, 26, 25, 1, -12, 14, 11, 6, -8, -4, -12, 12, 32, -8, 0, 16, 12, -2, -9, -9, -33, 5, -28, 6, 4, 7, 4, 18, -2, 0, -20, -48, -35, -16, -18, -14, -5, 11, -17, 3, 36, 37, 18, 7, 15, 12, -19, -43, 6, 29, 6, 3, 6, -7, -5, -10, -8, -22, -38, -51, -61, -63, -50, -39, -26, -52, -27, -14, 26, 12, 7, 11, 4, 9, -1, 5, 10, -51, -55, -35, 14, 20, 42, 43, 50, 32, 32, 33, -8, -13, -45, -46, -59, -81, -36, -3, 20, -17, -63, 3, 10, 19, 8, 9, -34, -44, -61, -42, -16, 19, 11, 29, 53, 29, 61, 50, 81, 55, -17, -28, -54, -54, -24, -42, -11, -19, -19, 0, 0, -6, 13, -20, -38, -50, -27, -35, -33, -10, 15, 24, 34, 11, 9, -14, 7, -10, -1, 1, -43, -12, -22, -82, -72, 7, 21, 11, 17, 10, -14, -2, -4, -2, -11, -19, 0, 7, -12, 19, -9, 31, 14, -5, 14, -8, -22, -12, -11, 0, -36, -31, -25, -39, -3, -3, 18, 16, -17, 0, 8, 42, -35, -20, -12, -34, -19, -32, -23, -34, -27, -17, -6, 9, 4, 47, 10, 10, -4, 3, -20, -20, 4, -10, 14, 9, -14, 4, -9, 10, -10, -70, -21, -14, -47, -23, -44, -45, -93, -56, -23, 40, 1, 0, -4, 28, 11, 20, -4, 16, -20, -9, 3, -12, -4, 3, 6, -44, -1, -42, -34, -27, 9, -6, -19, -18, -20, -48, -2, 2, 11, -18, -3, 24, 39, 32, 22, 64, -1, 1, -8, -17, -3, -31, -13, -31, -24, 18, 23, -16, 10, 1, -5, 3, 16, -6, -21, -16, 13, 7, 31, 36, 35, 26, 22, 44, 3, 18, -14, -20, 5, -27, -42, -54, -45, -11, 16, 17, -9, -4, -4, 6, 2, 21, 7, 9, 22, 30, 14, 24, 40, 11, 14, -1, -33, -1, -11, 2, 13, -13, -31, -50, -18, -19, 8, -26, 21, 26, -3, 11, 2, -17, 10, -12, -8, 1, -9, 43, 58, 30, 33, 45, -8, 7, -7, 3, -3, -56, -34, -42, 14, -28, -16, -26, 17, 7, 11, 15, 3, 11, 9, 15, -5, 5, -6, 20, 33, 7, 7, 38, 20, 0, -16, -18, 0, 14, -32, -20, -13, -11, -30, -17, -17, -18, -40, -31, -8, 0, -5, 5, -4, -11, -38, -32, -37, -24, 32, 79, 29, 16, -11, -5, 10, 16, -5, -28, -49, -48, -36, -56, 3, -9, -35, -3, -33, -25, -38, -3, -13, -34, -16, -25, -28, 21, 30, 33, -10, 4, 14, -14, -18, 2, -5, -30, -38, -1, 12, -23, -21, -54, -28, -21, -60, -27, -40, -25, -43, -32, -42, -7, 0, 1, -13, -30, 9),
  43 => (-12, 17, -13, -15, 13, 0, -13, 0, 13, -1, -4, -15, 4, 11, -10, 3, -33, -14, 1, 7, 5, -13, -19, 14, -4, 3, -12, 12, 8, -3, -17, -7, 16, -7, 6, 13, -9, 0, -6, 40, -11, 1, -30, -46, -54, -47, -46, -35, 3, 17, 12, -19, 4, 1, -12, 4, 19, -17, 20, -11, 8, 5, -9, 20, 17, -1, 52, 3, 26, -34, -40, -17, 1, -2, 36, 18, 23, 43, 15, -20, 26, -19, -18, -10, 10, 16, 19, 21, -12, 16, -10, 19, 35, 62, 85, 76, 7, -15, -8, 5, -24, 17, 33, 38, 2, -38, 28, -21, -15, -2, -7, -2, 8, 9, 17, 18, 8, -1, -18, 27, 4, 45, 50, 28, 12, -11, -8, 18, 8, 32, 20, 25, -22, -43, -4, 4, 4, 7, 6, -14, 10, -18, -1, 18, 2, 8, 22, 50, -37, -21, -33, 24, 22, -8, -4, 5, -8, -2, 11, 9, -51, -18, 9, 2, 8, -7, 13, -20, 13, 20, 1, -8, -13, -20, 32, 42, -29, 0, 19, 28, 14, 13, -8, 9, 20, 34, 10, -9, -14, -28, -32, -28, -4, -25, 25, 2, 10, 20, 16, -8, -13, -11, 51, 9, -12, 20, 3, 1, -16, 20, -4, 5, 36, 59, 41, -39, -42, -31, -46, -6, -18, -27, -7, -18, 13, 0, 16, 11, 6, 15, 37, -20, 3, -28, -10, 17, 13, 11, -9, 5, 12, 12, 2, -68, -53, -30, -60, -8, -21, -9, 3, -3, -19, 9, 2, 1, 8, -13, 16, -52, -75, -67, -41, -11, 17, 26, 8, 7, 19, 22, -47, -68, -15, -39, -63, -6, -35, -48, -47, -26, 15, -5, -15, 14, -7, -2, -51, -97, -83, -87, -7, 18, 38, 1, 1, 18, -3, -27, -51, -51, -18, -46, -44, -4, -29, -18, -10, 23, 17, 0, 19, 15, 6, -27, -82, -132, -56, -40, -4, 19, 39, 10, -4, 24, -17, -41, -33, -40, -17, -25, -22, 11, -16, -29, -2, -17, 12, -7, 3, 1, -3, -21, -115, -90, -25, -45, -5, 5, 55, 62, 30, -10, -33, -28, -55, -28, -16, -43, -17, 18, -34, -38, 7, -4, 5, -5, 11, -8, 13, -6, -42, -31, -39, 22, 56, 72, 84, 44, 19, -10, -44, -54, -26, -19, -6, -5, 42, 23, -22, -30, 5, -10, -7, 0, 17, -4, 16, 39, 1, 2, 6, 15, 43, 65, 45, 13, -6, -59, -43, -49, -30, -23, -53, -15, 36, 19, -13, -2, 3, -17, 11, 3, 16, -5, 14, 29, -23, 35, 47, 40, 46, 35, 9, 37, -17, -46, -13, -27, -23, -38, -23, -10, 12, -23, -8, 20, 6, -19, -16, -10, 2, -3, 3, 5, 9, 40, 48, 27, 44, 32, -20, -4, -44, -17, -35, -37, -2, -18, -32, -11, -12, -44, 13, 8, -12, 19, -7, -2, 6, -3, 39, -25, 24, 38, 11, 54, 78, 16, -2, -28, -50, -47, -44, -27, -4, -26, -29, -47, -43, -46, 28, 15, -19, -13, 1, 8, 8, -18, 3, -36, -8, 41, 17, 57, 40, 3, 11, -7, -7, -31, -40, -27, -25, -45, 0, -32, -13, -49, -4, 6, -19, -1, 13, 10, -5, 17, -8, -3, -14, 40, 32, 41, 27, -14, -6, 1, -24, -50, -47, -17, -37, -66, -34, -27, -13, -44, 14, 19, 24, 13, 2, 9, -13, 3, -20, -7, 34, 43, 15, 54, -7, -10, -26, -57, -44, -49, -46, -39, -50, -58, -16, 2, 11, -31, -3, 46, -1, 4, 8, 15, 2, 13, -29, -3, 58, 23, 42, 10, 14, -15, -11, -23, -34, -36, -53, -44, -47, -93, -4, 18, -8, -37, -43, -18, 3, 11, -1, 2, 2, 0, -61, 15, 68, 33, 15, 1, -19, -21, -20, -7, -45, -24, -39, -18, 2, -40, -39, 13, 0, -34, -24, 0, -15, -12, 12, -16, -3, -6, -16, 5, 28, 14, 18, -8, -19, -41, -25, -15, -28, -1, -11, -14, -19, -44, -24, 14, 31, -12, 7, -14, -9, -15, 9, -16, -18, -5, 34, 14, 33, 21, -14, -13, -13, -7, -24, -13, -21, -3, -14, 2, -11, 0, 3, 12, 1, -16, 14, -15, -4, 4, -12, -14, -2, 17, 6, 31, 50, -9, -31, -41, -32, -25, -24, -13, -19, -7, 12, -19, -2, 16, 14, 23, 32, 54, -16, 8, 7, 15, 15, -7, -14, 13, 2, 48, 27, 22, 6, -51, -53, -59, -45, -49, -3, 3, 26, -30, -4, -8, 23, -25, 21, 22, -25, -3, -9, -18, -8, -4, 1, -15, 6, 29, 38, 6, -3, 0, -52, -34, 3, -40, -32, 4, 18, -12, -31, -14, -21, 22, -24, 13, 0, -14, 13, 9),
  44 => (13, 1, -7, -6, 10, -5, -9, 10, 2, 0, -6, -17, -14, -17, -6, -63, -81, -34, -46, -55, -46, -65, -15, 20, 15, 17, -19, 1, -4, -15, 17, -6, 10, -17, 3, -11, -11, -20, 48, 48, 39, 18, 21, -21, 13, 14, 18, 24, 0, 23, 43, 26, 5, -10, 10, -17, 17, 20, -10, -6, -20, -9, 20, -12, 1, 51, 46, 74, 33, 1, 27, 8, 7, 12, 65, 51, 52, 9, 13, -6, -26, -18, 0, 16, -4, 2, -16, -6, 4, -21, 10, 18, 61, 73, 87, 51, 44, 53, 31, -3, 9, -25, 23, 27, 27, 41, 22, -19, -15, -28, -13, -10, 18, -2, -17, 16, -13, 6, 10, 43, 75, 70, 47, 62, 45, -15, -17, -14, -17, -35, -23, -13, 7, 30, 64, 1, -13, -4, 6, 15, 20, -7, -16, 5, -12, 1, 31, 46, 28, 61, 68, 69, 47, 27, 0, 3, -18, -24, -14, -14, 5, 7, 9, 32, -13, -35, -2, 11, 9, 17, 19, 7, 3, -6, 27, 89, 57, 77, 45, 61, 35, 41, 11, -15, -23, -32, 16, 8, 11, 36, 17, -9, 8, 1, -3, 11, -1, 9, 18, 3, 10, -13, 59, 85, 86, 54, 18, 13, 25, 35, 21, 26, 3, -25, 7, -4, -19, 39, 18, 13, 53, 7, -13, -7, 17, -6, 17, -17, 14, 18, 35, 63, 60, -5, -35, -14, 18, 45, 33, 32, 29, 34, 24, 20, 19, 34, 36, 34, 60, 8, -4, 7, -7, -8, -11, 2, -4, 1, 27, 42, 21, -5, 16, 15, 15, 48, 33, 35, 7, 17, 22, 17, 3, 26, 23, 45, 17, 29, 1, -15, -8, -9, 9, -2, -20, -16, 21, -7, -18, -13, -12, -29, 8, 30, 21, 40, 29, 23, 2, -3, 9, -4, -4, 34, 22, 5, 7, -19, -11, -14, -12, 20, -16, -29, -32, -85, -37, -43, -20, -35, -14, -17, -2, 62, 24, 9, -14, 19, 11, 5, 12, 8, -49, -20, -21, -13, 15, 16, -5, 13, -6, -26, -35, -69, -49, -48, -37, -23, 3, -8, 42, 64, 38, 16, 17, 22, 33, 9, 13, -13, -7, -31, -15, 13, 14, 7, 7, 9, 31, -24, -33, -59, -23, -29, -39, 5, 25, 9, 26, 88, 78, 32, 41, 34, 36, -16, -6, 9, -11, -26, -50, -29, 3, 17, 5, 18, -8, 24, -31, -5, 13, -9, -37, -10, 34, 31, 41, 43, 55, 29, 22, 27, 20, 3, -19, 22, 20, -1, -28, -14, -19, -8, 10, -16, -1, 17, -24, 15, 44, 1, -4, -4, 20, 79, 55, 40, 57, 20, -3, 55, 2, -9, 22, 23, 36, -7, -22, 21, -14, -8, -19, -7, -3, 27, 32, 62, 53, 16, 44, 39, 89, 73, 72, 47, 36, 6, 8, 30, 16, 6, 19, 53, 19, 8, -36, 37, 20, -9, 11, -2, 37, 58, 62, 58, 52, 19, 44, 18, 35, 64, 54, 41, 62, -9, 9, -7, 42, 36, -2, 17, 18, 15, -53, -4, -7, 3, 3, 18, 33, 38, 49, 51, 49, 41, 19, -1, 10, 9, 6, 19, 13, -3, -2, 15, 24, 12, 21, 14, 12, -29, -46, -41, 18, -7, -8, -15, 54, 30, 65, 37, 45, 5, -34, 9, -3, 6, 21, 34, 59, 34, 9, 23, -12, -13, 16, 54, 25, 20, -19, -50, 12, 14, -13, 6, 61, 66, 52, 1, -13, -24, -26, 21, 29, 14, 36, 18, 10, 36, 19, -1, 20, 1, 50, 55, 29, 2, -24, -38, 8, -13, -8, -10, 35, 48, 68, 51, 31, -9, 15, 18, 58, 40, 50, 44, 23, 32, 11, 55, 43, 44, 37, 41, 51, 50, 0, -4, 6, -4, 18, -13, 61, 62, 59, 28, 11, 4, 17, 10, 24, 37, 67, 65, 42, 54, 30, 52, 23, 29, 32, 53, 41, 8, 25, 53, -5, 4, 19, -16, 25, 44, 25, 19, 40, 3, 8, 24, 2, 22, 24, 26, 57, 43, 35, 31, 44, 59, 32, 17, 43, -2, -8, 43, -11, 18, -19, 2, -2, 44, 31, 41, 1, 21, 20, 58, 30, 44, 36, 55, 61, 45, 67, 31, 75, 66, 5, 14, 3, -15, 7, -19, 0, 7, 9, 3, -1, 24, 31, -11, -7, -11, -15, 19, 8, 27, 33, 40, 22, 32, 23, 32, 27, 47, 35, 13, 21, 1, -6, -33, 17, -11, -6, -12, 3, 11, 35, 23, -19, 6, -14, -4, -28, 23, 12, 28, 37, 9, 4, -22, 9, -10, 32, 27, 16, -14, -50, -34, 12, 16, 9, 6, 13, 48, 52, 69, 81, 41, 7, 20, -5, 3, -3, 22, 4, 25, 12, -16, -6, -26, -13, -5, 28, -7, -43, -25),
  45 => (16, -7, -11, 14, 10, 0, -16, 19, 16, 17, 15, 20, -20, 0, 28, -5, 7, 39, -7, -40, -23, 27, 10, 8, 7, 5, -20, 14, 17, -17, -10, -8, -16, -5, -9, 20, 1, 13, 10, -12, -8, 13, 44, 79, 68, 53, 52, 26, 17, 24, 53, -19, -30, -10, -8, 15, -18, 9, 15, -4, -15, -20, 20, 0, -3, 0, 1, 6, 80, 100, 69, 89, 33, 28, 22, -18, 9, 19, 11, -21, -42, 10, -15, 15, 6, -19, 5, -12, 16, 20, -3, 8, 2, -25, -14, 36, 30, 49, 43, 3, 25, 34, 20, -7, 6, 3, 43, -4, -6, 12, -2, -7, -17, 1, -12, -18, 13, -9, -17, -13, -48, -42, 22, 25, 4, 22, 12, 11, 32, -15, 13, -23, -19, 38, 30, 5, 12, 3, -7, -14, -13, 18, 4, -19, 4, 3, 3, -50, -24, 12, 7, -26, 8, -3, 31, 21, -3, -28, -13, -16, -39, 21, 8, 48, 17, 10, 0, 10, -8, 1, 12, -16, 20, 11, -33, -9, -14, 15, 31, -11, 17, 26, 28, -10, 9, 22, 29, 21, 28, 28, 40, 65, 33, -5, -17, -12, 11, -13, -17, -6, 9, 8, -37, 6, -2, 45, 29, 22, 33, 35, 35, 32, 6, -10, 33, 54, 12, 41, 42, 23, 0, -11, 51, 16, 18, 4, 14, -10, -11, 9, 8, 57, 46, 55, 24, -21, 14, 33, 43, 76, 15, 15, 40, 31, 2, 26, 31, 26, 22, 52, 35, 20, -3, 4, 12, -7, 12, 18, 31, 17, 22, 30, 23, 22, 25, 35, 45, 72, -1, 26, 37, 19, 38, 22, -9, 13, 10, 63, 44, 41, -11, 2, -8, 19, -6, -6, 52, 66, 69, 33, 16, 30, -7, -17, 16, 34, 19, 37, 22, 22, 36, 45, 13, -28, -29, 39, 53, 33, -2, 5, 18, -5, -2, -43, 65, 101, 88, 57, 32, 9, 7, 30, 17, 42, 28, 40, 21, 10, 53, 33, -1, 2, -6, -1, 29, 4, 7, -13, 19, 0, 4, -25, 67, 88, 105, 118, 77, 47, 72, 65, 91, 91, 69, 44, 31, 14, 48, 37, 22, 24, 6, 9, 4, 13, 11, -16, 10, -5, -40, -24, 37, 76, 96, 86, 65, 79, 65, 84, 85, 69, 86, 91, 54, 39, 72, 36, 75, 32, 69, 38, 41, 18, -1, 21, -18, -20, -33, -7, 66, 54, 47, 37, 48, 22, 32, 17, 18, 69, 84, 49, 37, 49, 50, 44, 76, 50, 63, 38, 31, -14, 2, 14, -2, 15, -16, 10, 67, 79, 41, 31, 47, 11, 30, 16, -25, 9, 20, 34, 19, 4, 2, 28, 44, 79, 58, 20, 40, 1, 3, -18, 10, 6, 10, 29, 52, 15, 40, -5, 39, 52, 4, -6, -20, 3, 10, 27, 23, -6, 21, 35, 19, 51, 22, 13, 29, -10, 9, 5, -17, 3, -2, 40, 30, 11, 9, 32, 15, -3, 16, 12, 29, 20, 33, -11, 14, 6, 7, 26, -3, 26, 7, 24, 35, 19, -13, -1, 8, -3, -16, -16, 15, 27, 10, 18, 18, 18, 36, 20, -4, 13, 26, 8, 22, 15, 5, 7, -6, 15, -4, 37, 41, 13, 15, 4, 20, -18, 5, 13, 26, -5, 44, 37, 13, 34, 9, 21, 14, 23, 14, 23, 24, 6, 18, 8, 11, -26, 4, 27, 24, 15, -11, 6, 13, -16, -19, 7, 70, 36, 37, -8, -7, -6, 0, 5, 5, 8, -6, -9, -9, 5, 34, -24, 14, -57, -19, 11, -11, -10, -5, 15, 20, 15, -13, 27, 25, 8, -12, 9, 8, -21, 10, 29, 15, 20, 7, 15, 4, 17, 19, -14, -11, -38, 12, 18, -47, -47, 9, -14, -10, 12, -34, -5, 7, 9, 3, -24, 10, -18, -16, -5, -10, -16, -23, -37, 13, 38, 18, -16, 8, -7, 26, -12, -64, -73, 2, 20, -5, -16, -26, -28, -27, -6, -34, -14, -27, -29, -3, -4, -28, -30, -21, -13, -14, 8, 19, -21, -13, -22, 4, 13, -17, -53, 20, -7, -7, -13, -28, -55, -49, 1, -32, -5, 19, -9, -18, -12, 0, -12, -48, -48, -25, -19, -46, -30, -30, -8, -12, 4, -26, -52, 0, 16, 0, 17, 0, -8, 37, -14, -2, 14, 30, 35, 6, -19, -24, -21, -13, 13, -24, -14, -28, -49, -68, -37, 10, 23, -49, -89, 3, 11, 10, 13, -37, 33, 17, -25, 12, 9, 40, 2, 13, 12, -4, 13, 23, 37, 29, 30, -10, 25, 2, -15, -10, 16, -40, -62, 19, -11, 1, 7, -15, 23, 47, 72, 62, 53, 84, 65, 56, 36, 17, 19, 32, 82, 67, 5, 28, -24, -28, -45, 24, 14, -41, -19),
  46 => (-11, -6, -7, 2, 15, -4, -17, 7, 19, 0, 4, 8, 14, 10, 3, 5, 18, 10, -26, -25, -37, -33, 12, 17, -17, -11, 16, -4, 18, 17, 16, -10, 15, 5, 17, -19, -14, 19, -21, -25, -18, -29, -34, -12, 8, 28, -22, -11, -25, -7, -36, -5, 2, 13, -11, -7, 18, 4, -13, -8, -5, -10, -3, -8, -17, -23, -28, -24, -45, 9, 34, 13, -33, -17, -24, -11, -38, -26, 3, -28, -6, 41, -18, 13, 10, 6, -17, 16, 7, -14, -9, 13, 5, 10, 61, 49, 29, 39, 0, 2, -8, -41, -8, 4, 2, -24, -31, 12, 5, -22, 0, -19, 3, 17, -6, 6, 8, 9, -2, -22, -11, 23, 29, 63, 46, 46, -17, -2, -2, -10, -17, -6, 1, -20, -7, 16, -6, 13, 6, -13, 11, -17, -14, -14, 11, -14, 6, 25, 16, 28, 50, 25, 2, -16, -23, -46, -28, 10, 5, -24, -15, 5, 15, 34, 34, 44, 0, 12, 3, 14, 13, -7, -11, 1, 36, 47, 37, 39, 30, -9, 26, 2, -28, -53, -6, -5, -9, 19, 13, 40, 19, -10, 5, -35, -16, 19, -7, 0, -5, 10, 1, -15, 21, 9, 31, 51, 20, -20, -21, -3, -56, -46, -8, 27, 23, 24, 29, 39, 15, 25, 22, 2, 1, -6, 4, 7, -1, -14, -7, -16, 0, 20, 51, 46, 10, -27, -13, -29, -35, -73, -48, 15, 27, 41, 65, 12, 18, 44, 20, 10, 0, 2, -9, 18, -6, 15, -20, -17, 39, 39, 70, 43, 27, -18, 3, -43, -80, -100, -22, 19, 22, 12, 23, 9, -3, 23, 40, 7, -21, 9, -19, -20, -4, -19, 2, -14, 32, 66, 53, 45, 9, -31, -34, -66, -44, -51, -22, -1, 11, -33, 1, -1, 13, 31, 33, 35, -34, -13, -4, -8, -11, 15, -14, 25, 21, 51, -1, -7, -10, -9, -28, -45, -49, -66, -24, 7, 31, 20, -7, -17, 8, 54, 32, 36, -3, -25, -18, 1, 20, -20, -19, -2, 27, -4, 17, -12, -10, -18, -37, -77, -63, -63, -63, -3, 4, 20, -23, -10, 5, 39, -9, 2, -33, 15, -18, 20, 7, -19, -15, -6, -1, -37, -5, 22, -32, -65, -92, -106, -100, -44, -70, -25, 8, 29, 20, -3, 31, 33, 28, -14, -23, 28, 17, 10, -4, -15, -10, 41, -7, 0, 33, 1, -20, -80, -88, -110, -65, -63, -73, -15, -22, 26, 32, 30, 24, 7, -16, -23, -56, 4, -8, 10, 13, 17, -4, 43, -4, -2, 55, 19, -17, -88, -84, -30, -36, -32, -48, 7, 35, 53, 58, 16, 20, -3, -1, -10, -19, 23, -14, -1, -18, -12, 3, 59, 24, 0, 67, 45, -5, -34, -45, -7, 13, -42, -55, 4, 54, 16, 78, 11, 29, -14, 12, -3, -32, 1, 19, 14, 17, 10, -11, 23, 18, 35, 57, 0, -30, -14, -27, 36, 1, -21, -8, 26, 58, 46, 36, 10, 16, -1, -9, 6, -10, 15, 16, -5, 4, -17, 25, 37, -12, 23, 24, -38, -55, -19, -6, 32, 26, 4, 5, 18, 12, 7, 35, 42, 21, -15, 4, 9, 4, 5, 17, 8, -17, -16, 23, 32, 0, 39, 19, -76, -102, -35, 22, 14, 23, 37, 9, 16, 43, 13, 26, 6, 29, -34, 5, 16, 4, 28, 6, -17, -11, -19, 23, 16, 44, 47, 6, -63, -31, -15, 10, 21, 24, 27, 30, 21, 48, 49, 9, 4, 38, -5, -12, 18, -55, 13, 11, 8, -10, -17, 22, 15, 14, 70, 6, -48, -19, 2, -24, 4, 42, -2, 23, 39, 50, 43, 48, 31, 8, 8, 31, 31, -37, 36, 1, 17, 9, 8, 42, -21, 27, 28, -13, -23, -12, -26, -24, -8, 29, 34, 29, 7, 27, 44, 32, 27, 12, -36, -5, 7, 11, 49, -17, -1, -7, 8, 18, 11, 3, -2, -35, -23, -48, -48, -3, -13, 34, 36, 44, 24, 29, 16, 18, 25, -30, -16, 5, 17, -45, 51, 18, -4, 6, 16, -6, -34, -24, 2, -7, -6, -19, 5, -4, -24, 31, 55, 29, 16, -1, 0, -10, 6, -15, -15, 12, -4, -18, 49, -15, -9, -12, 17, 4, -18, -9, 11, 18, -3, -13, -7, -17, 7, 18, 40, 14, 32, 12, -22, 12, 22, -24, -6, 27, -18, -8, 43, -11, 16, 5, -8, 5, 14, 11, 7, 28, 43, -14, -26, 0, 20, 45, 33, 26, 12, 8, 5, 23, 6, -21, -18, 2, 1, 30, -1, -11, 7, 6, -16, 13, -7, 11, -15, -43, 17, 8, -12, -12, -2, 26, 3, 13, -2, -22, -23, -37, -60, -71, -58, -20, -18, 57, 15),
  47 => (0, -16, 4, 5, -5, -12, -10, 4, 20, 0, -16, -6, 11, -4, 9, 6, -15, -12, -26, 6, -26, -7, 7, -15, -5, 12, -13, -12, -4, -10, -5, 13, 11, -13, -9, 3, -15, 10, 0, 8, -7, -11, -6, 2, 0, -2, -17, 1, -24, -18, -29, -26, 23, 5, 5, 19, 19, -7, -9, 9, -5, 11, 12, 6, 18, 10, 5, 9, 0, 27, 2, -3, -33, -65, -59, -76, -68, -11, -21, 40, 34, -7, 10, -4, 9, 15, -9, 12, 6, -2, -4, -3, 3, -20, -24, 13, 29, 12, -24, -4, -74, -65, -85, -77, -21, -4, 6, 72, 47, 35, -2, -8, 18, 5, -3, 6, 8, -6, 6, 14, -36, -52, -19, -31, -7, -26, -16, -27, -41, -49, -45, -54, -44, -14, -1, 62, 59, 0, 0, -18, -4, -15, 2, -13, 11, 18, -10, -24, -61, -48, 9, 14, -18, 12, -18, -5, 5, -23, -16, -7, -14, 2, 34, 26, 3, 10, -9, -9, -13, 13, 0, 13, -6, -16, 0, 11, -37, 12, 63, 71, 66, 44, 23, 12, 20, -18, -1, 5, 21, 2, 30, 22, 19, 33, 12, 3, -6, 16, -5, 15, 18, -16, -8, -20, -8, 46, 83, 55, 43, 36, 1, -24, -3, 19, 32, 48, -2, -11, 45, 40, 26, 15, -17, 2, -10, -15, -1, -9, -12, 14, 31, 15, 47, 45, 25, 66, 19, 34, -7, 1, -4, 7, -5, 36, 15, 33, 35, 40, 37, 10, 22, -46, 9, 2, 17, 13, 7, 20, 15, 28, 16, -38, -24, -42, -7, -8, -23, -3, -3, -22, 31, 28, 13, 18, 26, 15, 38, 8, -20, -25, 4, -14, -13, -7, -17, -35, 6, -56, -51, -109, -139, -124, -135, -93, -74, -15, -28, -12, 44, 44, 12, 43, 50, 28, 1, -20, -26, 2, 14, -9, 17, -3, 12, 0, -38, -102, -122, -128, -134, -101, -61, -83, -27, -16, -26, -28, 1, 27, 42, 51, 28, 22, -33, -18, -6, -32, 5, -1, 11, 6, -18, 22, -121, -138, -126, -79, -32, -17, -42, 21, 14, 18, 0, -11, 3, 4, 57, 20, 25, -12, -47, -27, -36, -25, -5, 11, -6, 5, 16, -34, -76, -99, -110, -29, -16, 13, -6, 18, 9, 13, -2, 5, 2, 13, 33, 19, -17, -21, -24, -22, -20, -7, -3, 6, 6, 15, 35, 24, -12, 2, -34, 38, 22, 6, 14, 17, 5, 20, -1, -14, 13, 24, 5, -2, 4, -41, -10, -21, -28, 27, -8, -17, 18, 5, 51, 71, 25, 58, 38, 56, 31, 30, -20, 37, 15, 21, 36, 22, 45, -21, 12, -16, -11, -37, -14, -3, -18, 17, 8, -20, 15, 5, 37, 77, 68, 60, 51, 12, 36, 8, -11, -14, 34, 8, 18, 17, 47, 6, 13, 4, 13, -14, -24, -26, -48, 8, -9, 15, -17, -19, 44, 37, 55, 34, -15, -16, -11, 1, -8, -24, 9, -3, 23, -27, -1, 1, -15, 6, 0, -27, -51, 1, -33, -5, 8, 4, 16, 5, 63, 35, 51, 53, 46, 29, 31, -2, -4, 24, 14, 49, -10, -12, -1, 5, -34, 13, 10, -3, -16, 12, -17, -1, -9, -17, 8, -3, 29, 37, 28, 49, 13, 14, 44, 12, 9, -4, 13, 17, 38, 27, -20, -19, -11, 18, 11, -4, -8, 13, -24, 22, 16, 11, -2, 17, 15, 25, 8, 0, -41, -18, -28, 24, 25, -14, -23, 10, 7, 13, 31, 10, -24, -22, -5, -12, -63, -39, -34, -14, -15, -1, -15, 12, -3, -16, 4, -28, -33, -24, -1, 62, 12, 10, 12, 8, 1, 9, 32, -10, -2, -21, -13, -43, -60, -44, -27, -21, -16, 7, 0, -13, -25, -22, 49, 16, -3, -21, 6, 44, 33, -7, 26, 35, 17, 47, 37, 17, 26, -15, -5, -42, -46, -46, -10, -19, -15, 20, -3, 4, -6, 39, 1, -8, 3, 8, -39, 19, 16, 29, 18, -13, 11, 28, 49, 24, -6, -23, 33, 0, -51, -55, -48, 13, 6, -8, -20, -15, -2, 26, 29, -5, -27, -19, -10, 0, -7, -35, -9, -12, -1, -44, 38, 15, 24, 12, 10, -37, -41, -55, -18, 4, -19, 1, 4, -5, 5, 30, -30, -41, -34, -26, -12, -21, -49, -29, -21, -48, -80, -58, -29, -21, 9, 7, 29, -28, -48, 3, 4, 4, -20, 14, -3, 13, 8, 6, -24, -39, -45, 6, 17, 17, -41, -41, -7, -18, -52, -28, -33, -12, -7, -10, 20, 6, -9, 21, -6, -8, 3, -15, -13, 10, -21, -4, 28, 10, -29, -11, -9, 13, 12, -40, -3, -7, -26, -65, -5, 0, -11, -22, 3, 19, 6, -1, 17, -1),
  48 => (-13, 8, 16, -8, 0, 16, -4, -7, 5, -4, -11, -5, 20, 17, 14, 1, -33, -22, -1, -5, 8, -30, -8, -17, 11, -4, -13, -19, 9, 19, 0, 0, 18, -16, -4, 19, -3, 6, -8, 14, 28, 17, 5, -17, -13, -25, -8, 15, 16, -9, -20, -2, 9, -19, -7, 5, -4, -6, -13, -16, 3, -4, 0, -15, 8, -28, 11, 8, 4, -24, 8, -13, -35, -7, -19, 3, 1, 36, 7, -29, 11, -8, 14, -10, 2, -10, -20, -18, -13, 7, 17, 10, -33, 6, -4, -16, -17, -33, -30, -5, 0, 5, -4, 9, 0, 55, 69, 3, 4, -19, -1, -3, 12, 8, -6, -17, -19, -1, 4, 2, -22, -9, -46, -37, -58, -41, -26, 9, -3, -20, 1, -17, -12, 20, 90, 50, -11, 26, -1, -3, 18, -15, -16, -18, -11, -8, -14, -10, -11, 0, 18, -32, -14, 6, 3, -5, 1, -25, -17, 15, 23, -10, 41, 27, -9, 23, 13, -19, 18, 1, 17, -5, -5, 7, 8, -36, 7, 51, 23, 30, 10, 14, 23, 19, 22, -26, -19, -9, -29, -43, -21, -2, -19, -6, -22, -15, -4, 11, -7, -6, -18, -19, -10, -11, 0, 15, 34, -8, 15, -7, 2, 20, 29, -11, -5, 3, -18, -37, -28, -32, -30, -15, 19, -6, -19, 8, 10, 7, -4, 1, 17, -28, -50, -40, -20, -32, -41, -47, -47, 11, 17, 18, 5, -14, -17, -29, -28, -72, -38, -38, 22, 10, -7, -3, 6, 4, -12, -5, -9, -32, -67, -36, -15, -47, -18, 10, -14, 3, 16, 9, 22, -60, -23, -13, -4, -8, -35, -68, 16, -21, 7, -10, -17, 17, -12, 29, -7, -41, -17, 24, 22, 28, 23, 33, 34, -13, -12, -18, -3, -6, -20, -12, 10, 25, 20, 10, -1, 1, 16, -13, -4, 3, -10, -22, -13, 2, 19, 30, 44, 13, 36, 24, 13, 2, 9, -6, -23, -5, -11, -21, -21, 22, 10, 19, 61, 19, -6, 7, -20, -17, 13, -3, 12, 2, 1, -24, -13, -23, -26, -23, -16, -43, -49, -16, -24, -11, -42, 3, 20, 21, 40, 33, 63, 6, -1, -8, -18, 3, 5, 12, 4, -46, -54, -82, -111, -88, -91, -60, -18, -42, -40, 3, 19, 27, 35, 44, 26, 26, 39, 63, 40, -22, 12, -5, -5, -10, 6, 3, -31, -58, -59, -107, -102, -86, -10, -9, 22, -20, 44, 43, 11, 43, -4, 14, 21, 27, 44, 11, 31, -39, 11, -19, -16, 6, -22, 3, -33, -42, -37, -66, -51, -15, 33, 51, 48, 7, 29, 19, 26, 16, 0, 9, 2, -16, 33, -6, -42, -57, 15, -16, 20, 20, 14, -29, 18, -2, -3, -10, 48, 36, 49, 46, 25, 33, 58, 55, 36, 1, -38, -10, -15, -15, -40, -44, -6, -19, -16, -13, -1, -12, 21, 9, 25, 55, 59, 75, 64, 60, 46, 60, 23, 23, -1, 39, 27, -23, -24, -41, -34, -34, -25, -57, -23, -1, -17, 20, 10, 14, 21, 69, 44, 54, 73, 47, 25, 29, 11, 5, -32, -71, -76, -20, -34, 16, -8, -10, -24, 0, -4, -21, -15, -48, -20, 7, -1, -6, 57, 46, 46, 11, 25, -8, -40, -83, -95, -84, -76, -74, -68, -78, -47, -17, 19, 36, 39, 15, 36, 10, -5, 1, -12, 21, -2, 0, 17, 8, -21, -22, 1, -39, -48, -54, -50, -31, -16, -26, -15, -33, 22, 1, 24, 15, 54, 46, 37, 13, 1, -15, -19, -6, 10, 8, 8, -40, -91, -65, -54, -39, -25, -44, -46, -21, 19, 49, 23, 9, 32, 5, 43, 25, 43, 41, 41, -50, -28, -19, 20, 1, -6, -19, -31, -16, -45, 4, -24, -53, -24, -38, 11, 27, 22, 35, 21, 35, 32, -9, 10, -5, 32, 28, 25, -42, -29, -41, -3, -8, 4, 4, -19, -13, 15, 21, 3, 37, 26, 21, 45, 31, 11, 7, -1, 32, 27, -9, 15, -5, 0, 12, -17, -57, -31, -30, 6, 4, 15, 2, 2, 31, 50, 53, 35, 40, 12, 19, -5, 25, -4, 7, 60, 60, 37, 40, 18, 10, -7, -24, -28, -18, -17, -4, 8, 17, 3, -13, -32, 24, 50, 23, 36, 2, 24, 23, 16, -7, 8, 1, 19, 34, 3, 9, 2, -9, -16, -73, -67, -61, -26, -12, -19, -12, 13, -10, 2, -4, 52, 10, -5, -10, -13, 16, 11, 56, 29, 21, 30, -10, -10, 16, -5, -23, -40, -50, -25, -22, -35, -33, 1, 6, 1, -7, 2, 33, 23, 28, -13, 16, -9, -2, -19, 18, 30, 19, -12, 8, -2, -16, -19, -20, -35, -44, -28, -56, -18, -23),
  49 => (14, 16, -18, -8, 7, -12, -19, 13, 8, 5, 13, 7, -3, 8, 13, -7, -24, -23, 5, 15, 5, 9, 9, 6, -10, -12, -7, -7, -16, 8, 3, -12, 20, 5, 14, -11, -19, -11, 1, -16, -18, -11, -26, -4, 20, -35, -6, 34, 26, -10, -16, -12, -9, 0, -13, 5, -6, -4, -8, 15, -16, -18, 0, 17, 14, -6, -13, -6, -43, -29, 7, 57, 26, -13, -15, -58, -35, -36, -18, -6, -20, -7, 15, -16, 2, -1, 17, -9, -10, 13, -11, -4, -25, -18, -35, -44, 39, 33, 45, 3, -1, 12, 0, -8, -31, -66, -34, -35, -15, -6, -13, -13, -20, -19, -20, -8, -1, 8, -4, -8, -10, -54, -103, -29, 12, 15, 5, -40, -37, -4, 10, -11, -55, -95, -53, -25, -11, 5, 12, 2, -16, 19, -7, -9, 2, -17, 5, -1, -10, -85, -63, -8, 37, 1, -75, -44, -11, -16, 7, 9, -39, -83, -79, -60, -41, -6, 16, 11, -7, 1, -2, 9, 12, -14, 10, -20, -53, -79, -11, 43, 5, -31, -88, -34, 10, 15, -13, -6, 1, -54, -83, -62, -35, -1, 1, -1, 6, -20, -9, -15, -15, -3, -12, -42, -30, -12, -5, 20, 7, 0, -25, -25, -22, -11, -5, 25, -18, -35, -60, -52, -6, -9, 2, 20, 1, 15, 12, 20, -13, 4, -3, -17, -62, -24, -2, 3, 3, -22, -57, -90, -25, 27, -7, 1, -3, -41, -28, -32, -40, -51, 6, 8, 17, 13, -10, 5, 10, -1, -19, -64, -37, -4, -11, -25, 23, -12, -94, -80, 10, 17, -6, 27, -26, -51, -45, -29, -82, -30, 13, -5, 15, -19, -14, 16, 0, 7, -50, -52, -38, 13, -1, 15, 34, 1, -119, -130, -22, 49, 24, 43, -21, -37, -80, -37, -30, -28, 4, 3, -11, -18, 6, -21, -10, -26, -8, -49, -48, -3, 35, 8, 34, -37, -96, -100, -19, 8, 14, 14, 37, -2, -40, -55, -13, -21, -25, 5, -5, -3, -15, -5, 4, -29, -6, -65, -57, -34, 14, -8, 2, -24, -67, -72, -37, -14, 13, 27, 28, -9, -49, -31, -20, 0, -6, 19, 6, -10, 18, -7, -34, 25, 6, -35, -52, 25, 16, 19, 38, 1, -64, -51, -18, -20, -4, 18, 42, -5, -30, -20, -33, -17, -18, -20, -16, -13, -8, 4, -33, 19, -5, -20, -39, 27, 2, 16, 44, 31, -49, -38, -38, -30, 2, 20, 35, 38, -24, 16, 57, 8, -24, 10, 18, -18, -19, -21, -3, -6, -16, -25, 3, 27, -8, 14, 46, 47, -27, -37, -50, -19, -4, 33, 49, 37, 6, 22, 70, 47, 19, 43, -15, 1, 16, -11, -38, -30, -64, -37, 41, 41, 63, 70, 42, 16, 10, -33, -41, -43, -7, 5, 51, 46, 22, 46, 61, 12, 19, 17, 9, 12, -3, -6, -38, -30, -53, -14, 36, 41, 54, 37, 29, 41, -3, -8, -18, -36, 4, -10, 43, 53, 12, 31, 53, -5, -11, 5, -15, -14, 13, -10, -12, 36, -1, 8, 25, 26, 26, 39, 23, 26, 6, -10, 16, -9, -22, -8, 6, -7, 6, 34, 33, 19, -3, 33, 14, -5, 8, -17, 25, 50, 62, 22, -15, -19, -1, 59, 35, 40, 3, -35, -16, -30, -34, 20, 26, 13, -18, 6, 39, 16, 8, 39, 1, -15, -14, -19, 40, 59, 11, 0, -42, -11, -19, 24, 31, 11, 16, -25, -22, -7, -6, -3, -3, 12, -16, -14, -4, 20, 49, 46, -20, -17, 9, 11, -11, -38, -47, -56, -16, -69, -9, 20, 33, 8, 17, -17, 4, -31, -9, -39, -13, -30, 18, -10, 9, 23, 41, 33, 18, -7, -5, 14, -2, -47, -9, -56, -54, -70, -43, 16, 16, 8, -21, -10, -23, -2, -8, -8, 2, -9, -2, 23, 20, -2, 44, 34, 13, 12, 11, 9, -8, -43, -62, -45, -66, -65, -53, -33, 41, -33, -12, 1, -41, -17, 3, -10, -3, -8, 3, 7, 41, 49, 41, 32, 10, 8, 15, 3, 1, 0, -38, -62, -52, -40, -34, -11, 20, 4, 5, 25, -22, -29, 2, -21, -8, 1, -2, 21, 48, 47, 43, 40, -14, -9, 20, 7, -4, -35, -32, -33, -25, -24, -33, -53, 6, -16, 4, 51, 44, 39, 14, -11, 26, 19, 29, 36, 67, 9, 5, -5, 11, -15, -17, -9, -16, -21, -19, -52, -32, -26, -47, -51, -93, -11, 9, 18, 28, 25, 36, 15, 4, -4, 15, 21, 22, 9, -30, -46, -15, 1, -5, 11, 6, 6, -7, 14, -15, -25, -1, -24, -43, -47, 0, 19, 8, -24, 12, 17, -9, 28, 10, 47, 29, -27, -46, -32),
  50 => (-12, 11, -10, -13, 20, -12, -19, 12, 13, 12, 13, -3, 9, 3, 20, 11, -20, -31, -38, 1, 22, 30, -8, -1, 16, -15, -2, -10, 14, 3, -17, 13, -13, 19, -11, -2, -18, -18, -16, -4, 55, 23, 2, -20, 3, -20, 16, -4, 16, 0, 12, 36, 5, -15, -6, -7, 11, 18, -2, -10, -8, 4, -7, 4, -17, 27, 8, 2, 10, 2, 21, 55, 20, 35, 11, -7, -22, -1, 30, 63, 37, 21, 9, 1, -7, -3, 15, -8, -11, 0, 3, -12, 39, 3, -6, 57, 58, 64, 44, 47, 42, 21, 11, -2, -20, -23, 19, -19, 46, -9, -12, -16, 12, -10, 12, -8, -13, -11, 5, -7, 20, -12, 13, 53, 9, 30, 28, 11, -10, 2, 15, -17, -26, 19, -19, 11, -15, 6, -10, -6, -14, -14, 15, -8, -1, -13, -13, 15, -7, -13, 38, 9, -19, 1, -5, 1, -41, -6, 11, -3, 19, 1, -8, 0, -54, 23, 2, -2, -9, -7, -2, -10, 5, 7, -13, -25, 7, -4, 12, -20, 21, 17, 20, -5, 10, 6, -38, -26, -7, -7, -1, -40, -42, 7, -14, -4, 16, 11, -18, -4, 5, 10, -4, -17, 36, 7, 21, -15, -15, 8, -1, 7, -9, -12, -38, -42, -13, 30, 6, -43, -33, 8, -1, -13, -15, -19, -20, 0, -19, -13, 17, 7, 11, 24, -12, 0, 4, 18, -19, -51, -26, -35, -18, -67, -42, 1, -29, -23, -33, -6, 11, 0, 14, -19, -8, -10, 9, -5, -25, -36, -27, -57, -32, -29, -30, 0, -23, -36, -49, -29, -37, -45, -24, -33, -33, -37, -45, -6, 13, 8, 9, -8, 7, -10, -7, -17, -34, -47, -56, -57, -65, -46, -47, -35, -34, -56, -42, -46, -20, -57, -44, -39, -57, -42, -59, -26, -18, 27, 11, -2, -2, -10, -14, -35, -39, -82, -20, -52, -41, -56, -32, 2, -32, -38, -1, -17, -14, -21, -22, -30, -39, -21, -56, -63, -19, -20, -11, -5, 0, 7, -6, -41, -30, -38, -13, 10, 6, -13, -29, 0, 0, -16, 27, 17, 16, 20, 6, 46, 0, 30, 13, -5, -3, -45, -8, 17, -5, -14, 20, 26, -37, 2, 5, -16, -16, -3, 1, 16, -2, -20, 5, 10, 21, 22, 29, 33, 14, 50, 18, 10, 25, -34, -17, -2, 0, 3, 34, 68, 39, 54, 83, 53, 28, 20, 38, 20, 7, -12, -21, 10, 31, -17, 14, 46, 38, 52, 74, 2, 32, 17, 6, -5, -9, 7, 4, 75, 40, 58, 78, 80, 25, 23, 22, 40, 24, 26, 29, 28, 4, -25, 38, 40, 36, 63, 42, 25, 38, 32, -20, -4, 10, -19, 33, 70, 21, 60, 40, 60, 55, 23, 36, 41, 44, 41, 25, 23, 23, 50, 26, 38, 58, 23, 60, 27, 40, 10, 14, -10, 10, -3, -13, 59, 42, 81, 45, 34, 16, 9, 27, 52, 23, 39, 31, 15, 36, 41, 43, 13, 31, 35, 33, 6, 21, 44, 19, 16, 3, 2, 3, 6, 37, 27, 33, 18, 39, 42, 50, 28, 28, 41, 41, 12, 28, 19, 53, 12, 16, 13, 25, 40, -20, 55, -5, -11, -14, 3, 29, 29, 31, -4, -5, -7, 20, 46, 18, 3, 26, 49, 64, 57, 33, 40, 53, 10, -3, 19, 1, -3, -3, 37, -20, 1, -20, 2, -21, 8, 45, 2, -21, -38, -18, 39, 7, -11, 24, 20, 30, 16, 50, 20, 25, 47, 20, 20, -2, -32, -33, 11, -4, 17, -14, -15, -26, -28, -12, -6, -38, -46, -65, -26, -45, -12, -35, -40, -2, 2, -2, -16, -41, -12, -16, 6, -14, -9, -28, -12, 15, -10, -9, 3, -25, -60, -22, -34, -45, -88, -87, -32, -64, -49, -59, -85, -68, -83, -51, -58, -91, -79, -66, -77, -67, 11, -26, -5, -3, -13, -10, 2, -29, -56, -46, -18, 5, -30, -59, -68, -56, -58, -88, -91, -46, -51, -60, -64, -71, -104, -67, -95, -69, -24, -37, -29, 5, -21, -13, -13, -9, -2, -27, 11, 35, 3, -7, -39, -45, -78, -85, -59, -36, -39, -18, -49, -58, -96, -77, -65, -109, -35, -12, -20, -11, 3, 15, -15, 20, 13, 14, 17, 16, 13, 21, -15, -39, -65, -67, -58, -17, -16, -8, -27, -55, -74, -71, -54, -28, -50, -31, -4, 4, 11, -15, -19, 30, -6, 24, -37, -61, 17, 22, -7, -27, -21, -54, -44, -21, -16, -28, -38, -32, -25, -37, -40, -8, 8, 2, -20, 17, -17, 20, 12, -9, 1, -29, 34, 3, -32, -7, -16, -21, -12, -37, -11, -4, -39, -9, -52, -63, -15, -52, -24, 11, 11, -9, 10),
  51 => (15, 4, 12, 16, -14, -15, -18, -17, -10, 13, -17, -7, 4, -3, 0, 22, 7, 8, 13, 15, 6, -20, 1, 3, -14, 1, -16, -20, 6, 0, -14, -18, 19, -9, -11, 1, 5, -11, 7, -16, -14, 23, -22, 0, -21, -37, -23, 4, -29, -5, -38, 24, -21, -14, -20, -4, 18, -1, 14, 19, 18, 10, 1, -5, 13, -42, -20, -13, -25, -30, -66, 20, 54, 51, 29, -13, -11, -45, -33, -33, 7, -23, -7, 15, -19, 13, 10, 19, 13, -3, 15, 14, -17, 35, 14, -44, -21, -44, -32, -17, 2, -23, -21, -10, -16, -48, -30, -6, -8, 6, 13, 7, -4, 8, -12, 14, -7, -19, -17, -24, 49, -5, -20, -55, -72, -10, 18, 18, -19, -23, 17, 8, 19, -42, -44, -18, 10, 7, -12, -13, -20, -19, 9, -1, -16, -1, 4, 41, 14, 0, -41, -94, 5, 16, 20, 2, -21, -31, 26, 45, 9, -39, -56, -91, -13, 1, -6, 15, 6, 19, -2, 11, 2, 15, 21, 51, 24, -18, -76, -49, -4, 14, 22, -37, -56, -57, 5, 48, 27, 13, -49, -68, -32, -6, 2, 19, -10, 2, 4, -9, -17, 4, 15, 13, -32, -30, -41, -28, 32, 21, 6, -23, -62, -30, 61, 50, -6, 5, -11, -47, -36, -14, 1, 5, -14, -20, -10, -1, 3, 7, -21, -22, -44, -62, -57, -29, -1, -1, 10, -18, -50, -38, 76, 79, 37, 21, -11, -31, 3, -17, 0, -23, 9, 14, 7, -18, 2, 20, -10, -51, -37, -89, -51, 15, 43, 27, -9, -11, -90, -84, 8, 63, 56, 33, 10, 21, 0, 9, 20, -33, 20, 1, -7, 10, -6, -14, -17, -21, -8, -30, 28, 3, 23, 21, 14, -32, -96, -113, -45, 59, 56, 43, 2, -2, 5, -21, 30, 8, 7, 5, -7, -16, -4, -27, 1, 26, 6, -14, -47, 5, 18, 26, 33, -20, -118, -95, -18, 71, 50, 10, 0, -4, -21, -32, 0, -1, -20, -20, 18, -5, -19, 3, 20, -3, -22, -36, -52, -14, 25, 27, 33, 27, -62, -91, -25, 25, 17, 2, -16, -28, -46, -22, -37, 34, -20, -4, 8, -19, -5, 40, 29, 3, -28, -23, -55, -4, 19, 24, 45, -5, -58, -47, -40, -35, -11, 32, -11, -21, -20, -19, -26, -7, 2, 13, 14, 13, 15, 62, 63, 3, -31, -31, -7, 22, 19, -3, 21, 42, -42, -56, -51, -49, -1, 25, -9, 18, 4, -57, -7, 15, -7, 14, 20, 2, 2, 37, 42, 3, 14, -8, -20, -3, 5, 8, 17, 34, -26, -33, -39, -21, -22, 7, 5, 21, -18, -45, -17, 23, 0, -13, -13, -20, 55, 39, 24, 12, -11, -26, -57, 15, -2, -3, 19, 43, -8, -43, -37, -58, -11, -2, -7, -3, -24, -16, 17, 65, -10, 1, -4, -15, 26, 33, 31, 0, -24, -22, 3, 26, 26, 3, 22, 19, 13, -36, -43, -50, 14, 50, 12, 8, -7, -51, 35, 28, -14, 11, 0, -8, -7, 76, 42, -14, -37, -24, -9, -3, 6, 24, 34, 10, 4, -18, -54, -13, -5, 29, 19, -17, -34, -32, -12, -13, 15, 1, -16, 11, 4, 28, 40, 3, -13, -20, 4, 21, 24, 31, 12, 8, 22, -22, -34, -56, -33, 23, 39, 3, -23, 5, -20, -26, -8, 18, -8, -4, -30, 38, 51, 3, -25, -23, -9, 30, 42, 29, 18, -4, 0, -3, -20, -13, 29, 8, 28, 41, 16, -23, -12, 21, 19, 18, 11, 13, -25, 59, 31, -10, -34, -41, -33, -2, 0, 15, 21, 4, -20, -33, -12, 11, -13, 15, -8, 11, 31, -15, 9, -44, -15, 3, -11, -2, 3, 48, 23, 39, -17, -21, -12, -2, 17, -8, 10, 5, -5, -48, -36, -23, 0, -21, -13, 30, 24, 33, 15, -46, 3, 14, 20, 15, -10, 65, 11, 39, 31, -20, -29, -9, -15, 23, -8, 3, -37, -44, -12, -20, -27, -51, -27, -6, 8, 16, -5, 0, -13, 6, -6, -11, -8, 7, -4, 15, 23, -28, -8, 1, -9, -26, 29, 38, -1, -29, -24, -44, -48, -41, -81, -14, 14, 46, 44, -17, -6, -18, 8, -8, -2, -25, -22, -4, 22, -25, -18, -13, -13, 0, 14, 13, 15, -3, -41, -20, -35, -39, -13, -33, -1, 30, 15, -6, -10, -12, -8, -19, -41, -32, -57, 25, 13, 13, -29, -30, -12, 12, -1, 4, 1, -20, -41, -23, -21, -22, -10, -59, -11, -13, -21, 8, 2, 0, -1, -10, -2, -5, -45, -53, -1, 0, -28, 1, -17, 21, -21, 10, 33, 31, 13, 26, 4, -7, -50, -76, -40, 13, 15, -8),
  52 => (14, 17, 9, -1, -20, -15, 14, -18, -13, 16, -6, 6, 20, 12, 3, 7, -1, -10, 1, -11, -11, -40, -12, 8, 9, 13, 12, 19, 14, 14, -17, 19, -5, 13, 11, 19, 9, -20, 6, 13, -21, -12, 4, -7, 16, -18, -22, -28, -8, -26, -12, 5, -18, 5, 19, 0, 5, 13, 15, 12, -12, 3, -13, -18, -5, 5, -6, -14, -28, -1, -31, -40, -27, -31, 4, 26, 12, 58, 47, 37, 7, 11, -13, -7, 18, 6, -4, -16, -16, -8, -2, -6, -17, 11, -19, -51, -40, -56, -68, -20, 4, 17, 17, 31, 29, 62, 45, 16, 55, 17, 9, 20, 13, 19, -19, -10, -12, 12, -6, -8, -1, -42, -34, -35, -20, -35, -36, 9, 1, -5, 13, 19, 20, 16, -15, -19, 18, 16, -5, -17, 14, 1, -17, -15, -20, 4, 8, 10, -15, -69, -44, -39, -29, -42, -7, 35, 11, -16, 1, 27, 10, -16, -37, -15, -30, 7, 1, -3, 18, 16, 9, -14, 9, -8, -1, 22, -47, -21, -38, -35, -31, -21, 25, 6, 5, -9, 5, 10, 17, 5, -8, -2, 9, 5, 0, 5, -4, 18, 11, -16, 0, 1, 7, -17, -84, -76, -84, -29, -29, -6, 23, 3, -2, 7, 5, 37, 11, 5, -2, 20, 40, 32, -16, -6, 15, -16, 8, -3, -9, -2, 13, -79, -63, -65, -90, -43, -1, 34, 15, 26, 22, -18, 0, 20, -15, 11, 20, 18, 27, 49, 9, -44, 9, -6, 13, 6, -7, -8, -25, -39, -53, -68, -85, -72, -29, 42, 48, 33, 13, -16, -2, 6, -39, -24, 7, 21, 51, 59, 15, -35, 19, 15, -9, 9, -18, 22, -32, -41, -22, 10, -72, -84, -1, 10, 72, 35, 27, -8, -5, -5, -24, -17, -14, 8, 15, 39, 56, 39, -7, -1, -7, -5, -10, -15, -45, -18, 21, -8, -47, -60, 15, 17, 32, 27, 22, -7, -20, -41, -36, -22, 1, -29, 19, 39, 75, 18, -13, 15, -1, 2, 14, -45, -43, 31, 14, -50, -17, -52, 20, 46, 49, 45, 32, -12, -40, -11, -31, -5, -24, -46, -35, 33, 27, -4, 0, -15, 13, 6, -7, -34, -5, 19, -19, -50, -37, -63, 6, 47, 53, 54, 39, -35, -63, -51, -14, 6, -6, 6, -17, -1, 39, -10, -15, 5, -4, 4, -10, -7, 44, 33, -54, -103, -86, -75, -17, 7, 9, 43, 19, -41, -73, -49, -11, -11, 17, -29, 8, 29, 55, 32, -1, -10, -10, 16, 3, -17, 25, 50, -40, -87, -93, -94, 3, 36, 28, 26, 14, -33, -44, -20, 11, 15, -3, -4, 15, 21, 28, 10, -1, -2, -18, -4, 34, -5, 19, 49, -45, -92, -133, -68, -19, 17, 16, 44, 20, -21, -56, -18, 1, 15, 6, 26, 22, -10, 18, 9, 6, -4, -9, 15, -24, 15, 60, 62, -20, -116, -126, -66, 8, 1, 10, 6, -7, -29, -83, -16, 3, -4, 4, 23, 40, -14, -22, -19, -14, -6, -1, -6, 13, 35, 61, 33, -43, -122, -126, -105, -1, 18, 8, -1, -7, -42, -65, -36, -11, -1, -20, 12, -4, 19, -21, -36, 11, -2, -19, -1, 0, 42, 41, 24, -80, -106, -122, -118, -5, 25, 38, 4, 18, -8, -29, -27, -39, -18, -20, -32, -24, -11, -4, -39, -10, 13, 13, -11, -20, -1, 66, 35, -11, -93, -133, -73, -27, 27, -2, 0, 20, -13, -36, -6, -19, -2, -27, -10, 3, 22, 12, -28, -11, 18, 7, 5, -41, -5, 27, 36, -38, -84, -78, -62, -55, -15, -6, -20, 20, -6, -15, 2, 6, -9, 4, -3, 30, 24, 12, -59, 10, 16, -9, -9, -22, 13, 28, 32, -26, -54, -58, -74, -57, -37, 6, -1, 0, -3, -28, -9, -12, -4, 8, 8, -10, -25, -39, -32, -13, -5, -11, -19, -17, -20, 43, 33, 1, -15, -32, -43, -40, -20, -18, -8, 10, 7, -3, -22, -7, 6, -27, 4, -28, -29, -42, -26, 10, -15, 11, -6, -3, -7, 10, 23, 30, 7, -13, -42, -59, -53, -16, -23, 15, 13, 0, -30, 32, 0, 8, 17, -5, -74, -63, -26, -8, 11, 9, 2, 13, 7, -1, 14, 17, 5, -13, -8, -39, -53, -28, 7, 5, -12, 15, 10, -7, -6, 18, -10, -31, -69, -47, -34, 7, -11, 9, -6, -20, -5, -2, 3, 0, -6, 5, -20, -1, -24, -23, 6, 1, 3, 6, 7, 18, -12, -45, -36, -49, -53, -33, -30, 12, -7, 7, -19, 7, 19, -8, 4, 2, -12, 13, -25, 5, -18, -31, -6, -26, -34, 16, 31, -3, -25, -27, -48, -53, -66, -36, -8),
  53 => (-12, 19, -17, 12, -1, -8, -3, -18, 3, -5, 3, 17, -17, 5, 7, -55, -48, -16, -52, -20, -4, 23, -21, -8, 0, 6, 7, -10, 16, -8, 1, 6, -9, -15, -11, 5, 16, -10, 13, 29, 7, -2, 6, -30, 17, 48, 25, 17, 21, 54, 60, 2, -44, -12, -10, 0, 17, -17, 19, -15, 2, 5, -16, 6, -12, 53, 19, 15, 50, 49, 68, 38, 20, 51, 28, 12, 26, 52, 4, 54, -23, 17, 7, -20, -19, 7, -17, -9, -5, 3, 14, 16, 9, 13, 18, 53, 75, 79, 61, 34, 2, -10, -17, -13, -15, -13, 3, -13, -23, -43, -14, 1, 14, 12, 6, 18, -16, 2, -10, 8, 27, 20, 69, 90, 48, 59, 24, 20, -16, -27, -22, -11, -21, 5, 26, -9, -33, -24, -17, 10, 10, 15, 8, -7, -10, -6, 42, 55, 3, 59, 34, 63, 4, 23, 5, -10, -30, -43, -10, -16, -33, -2, 25, 1, -38, -11, 19, 5, -15, -5, 0, 14, 13, -5, -2, 43, 19, 26, 48, 11, 10, 27, 31, -15, -20, -3, -51, -29, -21, -1, 25, 26, -1, 38, -7, 15, -20, 18, -17, 5, -3, 7, 27, 73, 26, 45, 19, 8, 50, 42, 42, 36, 19, -40, -26, 19, 7, 4, -1, 25, 20, 21, -7, 12, -12, 19, 16, -5, -6, -14, 51, 55, 30, 43, 33, 8, 35, 48, 35, 18, 22, 26, 24, 22, -7, 14, -28, 20, -2, 31, -24, 10, -15, 19, -17, 0, 10, -14, 22, 13, -35, -12, -9, -18, -14, -11, 4, 20, -4, 3, 4, 23, 3, 23, 48, 49, 13, 25, 21, 15, 11, 0, -2, 7, 6, -23, 1, -33, -39, -41, -60, -26, -19, -16, -8, 18, 5, 12, 10, 11, 22, 63, 39, 8, 20, 24, 36, -1, -13, -12, -5, -5, 7, -67, 0, -53, -7, -56, -72, -24, -12, -13, 19, 60, 8, 23, 18, 12, 22, 18, -2, 22, -10, -11, 19, -14, -1, 3, -5, 1, 35, 32, 73, 4, -7, -16, -37, 7, 39, 17, 40, 61, 19, 60, 52, 26, 31, 13, -3, 8, 9, 8, 47, 38, 6, 19, 7, -8, 54, 85, 103, 73, 48, 34, 44, 23, 22, 36, 65, 54, 78, 77, 64, 69, 31, 29, 15, 19, -13, 67, 31, 35, -18, 16, -13, -3, 44, 47, 66, 59, 70, 86, 80, 53, 68, 62, 50, 95, 65, 85, 64, 32, 25, 68, 24, 3, 56, 79, 36, 37, 12, -8, -12, 8, 2, 25, 36, 55, 67, 89, 98, 76, 57, 20, 25, 66, 33, 37, 34, 0, 4, 17, 40, 34, 43, 57, 24, 42, 2, 10, -11, -18, 21, 42, 54, 56, 69, 68, 70, 26, 30, 24, 29, 75, 60, 57, 49, 23, -5, 17, 39, 37, 17, 39, -14, 54, -15, 15, -9, -6, 21, 48, 54, 45, 41, 28, 2, 11, 9, 50, 62, 59, 60, 40, 29, 0, -2, 16, 10, 35, 40, 39, 2, 64, -9, 0, 9, 16, 18, 48, 32, 23, 5, 4, -18, 14, 7, 40, 49, 34, 17, 10, 44, 15, 5, 0, 25, -4, 10, -2, -10, 0, -1, -15, -10, 3, 44, 59, 37, 20, -5, 26, -1, 19, -12, 18, 29, 33, 39, 50, 33, 2, 3, -6, -13, 24, -28, -18, -11, -29, 11, -5, 3, -16, 7, 50, 68, 16, 15, -10, -33, 9, 15, 23, 12, 23, 39, 24, 32, -3, 28, 19, 1, 6, -16, 10, -37, -31, -12, -18, 12, -15, -37, 62, 61, 38, 10, 14, 25, 13, 41, 41, 29, 41, 27, -8, 7, 11, -7, 9, -7, 13, -4, 4, -40, -48, 5, 9, -6, -17, -13, 10, 50, 39, 28, -16, 44, 40, 13, 24, 25, 32, -15, 14, -14, -12, -34, -3, -2, 14, 28, 3, -2, -30, -8, 1, 5, 11, 2, 50, 30, 13, 6, -30, -3, 5, -22, -16, -23, -27, -19, 9, -22, -9, -3, 9, 16, -23, 41, 14, 7, -4, -12, 15, 11, -6, 13, 32, -4, -17, -45, -30, 2, 32, 25, 8, -1, 21, -17, -23, -12, -11, 28, 25, 0, 15, 31, 16, 41, -22, 15, -4, 4, 7, 15, 29, 58, -22, -27, -26, -13, -15, -39, -37, 16, 20, 9, 4, -20, 3, 35, 31, -14, 3, 69, 85, 5, -18, -18, 19, 6, -13, -14, 28, 10, -15, -14, 1, -35, -32, -24, -21, 21, 21, 35, 21, 17, -18, 31, 27, 20, -24, 16, 45, -1, -8, -20, -2, 15, 0, 16, 27, 37, 75, 47, 5, 3, 18, 0, 4, 57, 39, 38, 60, 45, 3, -21, -15, -21, -8, 7, 3, -30, -8),
  54 => (16, -17, -19, 20, -14, 19, 5, -7, -12, 1, -11, -21, 20, 16, -18, 19, 12, -26, -17, -9, -36, -6, 13, -8, 8, -4, 9, 8, -13, -10, 13, 15, 20, 1, 15, 19, -17, -16, 8, 5, -46, -26, -1, -26, 4, -35, -38, -5, -26, -17, -9, 2, -9, -5, 14, -16, 15, -5, -14, -18, 7, 19, -19, -12, -2, 11, 2, -86, -15, 2, -11, -14, 28, 11, -6, -17, -2, 31, 2, -7, -29, -2, -14, 14, 20, 20, -11, 7, -1, 14, 19, 3, -21, -28, -66, -33, 11, 18, 21, 50, 49, 37, 2, 1, 9, 25, 7, 0, -21, 14, -7, 9, -9, -6, -11, -7, -2, 1, -16, -13, -38, 22, 29, 31, 60, 26, 11, 56, 45, 31, -3, 30, -6, -11, 42, 9, -15, 6, 16, -15, -7, 19, -5, 2, -4, -9, -11, -51, -22, 30, 29, 30, 16, 0, 39, 43, 33, 53, 18, -9, -10, -39, 8, 38, 5, -18, -10, 20, -13, 12, -19, 5, -9, -20, -28, -29, -7, 16, 27, -13, 46, 26, 38, 41, 39, 30, -7, -8, -21, -39, -6, 11, 10, -9, 29, -14, 20, -9, 20, 14, -6, 20, 6, 4, 19, 2, 0, 14, 10, -30, 15, 0, -7, 23, 30, 37, -14, -16, -14, -7, -12, 1, -3, -34, -6, 15, 10, 4, 11, 5, -27, 19, 19, -9, -16, 20, -52, -90, -77, -45, 2, 3, 30, 22, -47, -44, -48, -4, -21, -22, -15, -20, 9, -9, -8, -14, 18, -12, -38, -1, 0, -55, -45, -59, -102, -120, -80, -52, -27, -8, -9, 1, -10, -49, -25, 3, -18, 2, -21, -18, 11, -15, 17, -16, -8, 5, -57, -58, -46, -52, -73, -62, -36, -46, -20, -26, -13, -12, 18, -31, -48, -22, -24, -9, -21, -28, -19, -21, -1, -9, 19, -21, 12, -40, -55, -40, -33, -38, -4, -14, -7, 22, 29, 4, -7, 6, -18, -12, -12, 1, -11, -20, -6, -10, -17, -18, -15, 1, 3, -8, 20, -8, -37, 6, 40, 18, 46, 68, 9, 14, 32, 41, 22, -19, -33, 10, -23, -10, 17, -27, -36, -20, -23, -65, 14, 9, -6, 13, 8, 24, 12, 20, 18, 36, 42, 22, 11, 18, 29, 14, -6, -11, -36, -24, 7, -17, 13, 27, 9, 24, 15, -58, -4, -4, -8, -9, 54, 27, 41, 28, 36, -7, 20, -2, 16, -2, 40, 33, 32, -25, -7, -12, -21, -24, 15, 8, -4, 38, 16, 0, 16, -13, 11, 10, 58, 39, 33, -19, 8, -7, -10, 4, -9, -9, -19, 3, -1, -43, -59, -81, -58, -72, -36, -13, -30, 6, -7, 2, -8, -3, 5, -15, 31, 32, 14, -21, -27, -64, -65, -40, -40, -24, -28, -3, -31, -77, -78, -69, -61, -71, -22, 2, -10, -17, 1, 2, -17, 10, -5, -8, 23, -14, -4, -10, -18, -24, -43, -75, -46, -23, -46, 2, -13, -45, -46, -49, -52, -42, 1, 25, -27, -30, 13, -13, 13, -14, -5, 14, 9, -39, -45, 5, -21, -41, -53, -57, -35, 2, -20, -28, 3, -21, -45, -40, -40, -31, 4, 42, 1, -52, -4, 23, 9, -10, 14, 16, 12, -23, -22, -15, -12, -12, -31, -13, -35, 14, -6, -30, -23, -15, 9, -13, -29, -31, -13, -7, 5, -15, -11, 20, -20, 11, 2, -16, -17, -31, 1, 17, -31, -35, -51, 6, -27, -23, -20, -12, -27, 9, 24, 16, 24, 11, -5, 2, 7, -1, -20, 12, 15, 17, 5, -11, -15, -8, -24, -18, -38, -41, -12, -9, 1, -18, 6, 5, -8, -15, 27, 33, 47, 28, 55, 42, 8, 10, -5, 33, 1, 0, -19, -20, 7, -15, -4, -21, -11, 19, -11, -3, 30, -2, 35, 26, 19, 7, 24, 17, 49, 60, 54, 34, 13, 38, 26, 40, 15, 0, 16, 3, 4, 42, 41, 33, 22, 15, 19, 22, 10, 14, -7, 38, -7, 21, 10, 22, 8, 58, 45, 45, 7, 78, 73, 65, -17, -13, -15, 1, 27, 62, 32, 50, 45, 61, 13, 24, 12, 27, 31, 20, 32, 33, 27, 44, 53, 50, 54, 11, 20, 27, 30, 27, -6, -13, 4, -13, 30, 34, 88, 67, 32, 39, 28, 29, 17, 2, -27, -1, 12, 12, 36, 67, 41, 54, 52, 42, 9, 15, 23, -5, 19, 13, 5, 15, 19, 37, 35, 38, 34, 43, -9, 32, 25, -23, -17, -5, -10, 15, 47, 30, 28, 22, 28, 36, 11, -4, 34, 25, 7, 12, -8, -10, -2, 1, 5, 5, 25, 9, 31, -2, -30, -28, -15, 5, 0, -15, 34, 44, 36, 16, 30, 44, -14, -21, 21, 28),
  55 => (-3, 5, 14, -20, -7, -9, -20, 9, 2, 10, 9, 8, 14, 17, 5, -23, -5, -19, -35, -70, -26, -46, -8, -1, 6, -11, 9, -12, -21, -16, 20, 6, -14, -3, 20, -2, 3, -16, -10, -31, -24, -9, 17, 14, 8, -10, -46, -73, -60, -36, -34, 12, 18, 16, -19, 5, 16, 18, -16, 12, -6, -4, -20, -20, 7, -19, -17, -12, -11, 19, 18, -13, 8, -10, 14, 20, 28, -14, -11, 6, 42, 15, 10, -15, -2, -16, 1, -3, -20, 0, -20, -14, -33, -28, 9, -17, 11, -6, -1, 5, 7, 17, 58, 70, 25, 19, -47, 12, -6, -3, 20, 19, -13, -18, 2, 18, -5, -13, 18, -16, -17, -6, 1, 32, 32, -13, 19, 8, 15, 34, 23, 30, 38, -37, -64, -29, -24, 4, -9, -4, -5, -3, 14, 1, 6, 9, -32, 0, 10, -15, 31, 40, 22, 21, -39, 0, 12, 26, 29, 16, -16, -52, -48, -56, -19, 1, -19, 9, -10, -5, 17, 3, -8, 19, -21, -6, 25, 51, 32, 44, 33, -20, -34, -52, 11, 8, 0, 0, -40, -64, -67, -42, -40, 14, 12, -18, -14, 3, 3, -5, -2, -10, 38, -14, 57, 60, 20, 19, 44, -23, -74, -60, -34, 11, 6, 9, -6, -32, -46, -59, -39, 9, 0, -8, 17, 11, -12, 6, -18, -14, 5, 31, 106, 29, 29, 51, 50, 19, -40, -61, -47, 13, -23, -17, 38, 5, -31, -13, -37, -3, 9, 18, 20, 20, 16, 9, 2, -17, 30, 81, 84, 28, 39, 17, 43, -6, -48, -86, -32, 0, -9, -27, 36, -10, 14, 3, 42, -17, 2, -11, -21, 10, -16, -6, 9, 5, 65, 72, 70, 2, 2, -8, -2, -17, -46, -71, -20, 3, -22, 17, 19, 4, 8, 3, 31, 19, -27, 8, 9, 11, -3, -18, 21, -19, 11, 26, -10, 5, 1, 5, 26, -32, -36, -25, -9, -11, -15, 3, 33, -1, 14, 3, 23, -3, -9, 22, -3, -15, 18, 18, -8, -58, -50, -35, -51, -54, -6, -15, 9, -27, -52, -21, -27, -10, 18, 4, 17, -8, 0, 5, 12, 11, -10, 21, -12, 11, 5, -4, -55, -44, -33, -67, -74, -33, -18, -4, 16, -10, -9, 8, -43, 5, -5, -9, 16, -6, -34, -44, -3, -22, -4, -10, -7, 19, 19, 18, -36, -13, -81, -126, -67, -1, -30, -41, -15, 10, -1, -21, -43, 20, 21, 23, 18, -2, -45, -23, -30, -36, -36, -34, -11, 14, -4, -7, -9, -43, -104, -103, -78, -25, 17, 5, -16, 26, -21, -4, 5, 14, 18, -15, 7, -24, -39, -34, -31, -15, 24, 26, 2, 3, 16, 17, 15, -4, -37, -57, -32, -13, 1, 8, 34, 14, -7, -42, 4, 33, -13, 0, 25, 22, -31, -13, -49, -13, 25, 55, 9, -13, -6, -10, -7, -3, -76, -32, 25, -34, -5, -8, 20, 15, -15, -12, -37, 7, 20, 10, 9, 36, 6, 15, 0, 2, 35, 69, -3, -3, 13, -12, -6, -22, -30, -52, 2, 14, -22, 23, 34, -1, -4, -13, -19, 41, 35, 36, 36, 3, 27, -1, -39, -16, -8, 50, 0, 2, -9, -11, -12, -63, -44, -57, -20, 2, 20, -2, -4, -46, -60, -44, -44, 67, 43, 52, 47, 34, 10, -40, -29, -47, -12, 36, -12, 16, -9, 10, -12, -53, -41, -30, 20, 22, 0, 7, 13, -34, -54, -61, -33, 57, 58, 41, 42, 39, 2, -24, 3, -35, -21, 33, 18, 4, -8, -6, -8, -20, -29, -19, 13, 9, 41, 26, -48, -28, -89, -105, -91, 16, 39, 21, 0, 12, 0, -7, -34, -52, -22, 14, 6, 15, 1, 12, -32, -36, -47, 4, 12, 36, 44, -22, -75, -82, -110, -104, -76, 30, 57, 36, 43, 49, 36, 6, 12, -46, -45, -7, -18, -12, 3, 5, 5, 2, -29, 29, 38, 63, 60, -13, -38, -46, -90, -89, -70, -3, 49, 32, 51, 70, 57, 18, -9, -52, -56, -17, -1, -2, -9, -4, 1, 15, 25, 27, 21, 49, 43, -32, -45, -60, -57, -63, -31, 20, 16, 28, 9, 10, 28, -18, -18, -38, -40, -11, -1, -15, 0, 19, -8, 16, -27, 12, 14, 22, 28, 1, -65, -63, -81, -103, -30, 9, 48, 45, 36, 61, 58, -9, -37, -36, -20, -42, -13, -10, -10, -1, 21, -5, -13, 5, -30, -15, -7, -17, -28, -50, -81, -78, -78, -9, 41, 63, 54, 57, 30, 3, -13, -47, -41, -23, -6, -19, 8, 0, -8, 0, 10, 14, 11, -17, -39, -29, -25, -46, -54, -60, -36, -29, 5, 6, 6, 20, 22, -6, -10, -43, -41, -31),
  56 => (12, 4, 12, 16, 9, -10, -13, 19, 5, -16, -19, 0, 16, 4, -4, 0, -6, 13, 36, 18, 16, -6, 14, 20, -21, -20, 16, -5, -9, 0, 2, -16, 11, -3, -17, -6, -1, 7, -17, 4, 3, 12, -9, -10, -29, -11, -1, 20, 34, 22, 20, 23, -8, -14, 16, -10, 4, -5, 20, 15, 20, 7, -3, -8, -3, 16, -17, 6, -8, 1, -47, -58, -25, -11, 47, 21, 11, -3, -10, -6, 20, 19, -7, 11, 7, -4, 11, 16, -6, 19, -15, 17, -19, 18, -18, -19, -71, -86, -93, -34, 8, 20, -6, 2, -2, -11, -36, -6, 15, -20, 3, 13, 14, 17, 3, -2, 9, -4, -15, 9, 20, -22, -62, -67, -46, -54, -56, -29, 24, 31, 5, -3, -39, -37, -16, 13, -8, 15, -6, 18, -11, -15, -13, -7, -12, 6, 13, 10, -22, -46, -53, -94, -106, -57, -18, 29, 50, 64, 21, 2, -29, -28, -30, -12, -13, -35, 20, 8, 18, -8, -17, 2, -1, 1, -8, -51, 52, -1, -62, -103, -107, -86, -33, 33, 14, 72, 5, -29, -63, -44, -60, -69, -38, 0, -21, 9, -5, -17, 5, 0, 6, -11, -44, -51, 13, -42, -45, -70, -95, -82, -37, 44, 12, 18, -11, -66, -70, -41, -43, -43, -43, -14, -3, 14, -13, 3, 16, 13, -17, -9, -6, -32, -33, -10, -23, -47, -76, -99, -19, 3, 6, -6, -8, -22, -3, -8, -49, -50, -59, -45, 1, -5, 5, 7, -5, 2, -19, -11, -7, 13, -13, -23, -35, -36, -91, -74, -19, -21, -9, -32, -23, -39, -23, -24, -29, -71, -34, -35, -27, -8, 10, -3, 15, 0, -1, -10, -18, 13, -89, -35, -31, -48, -79, -68, -68, -27, -29, -26, -11, -12, -48, -15, -14, -45, -30, -16, -14, 2, -20, 14, 6, -7, 6, 19, 42, 15, -22, 12, -8, -25, -69, -56, -12, -10, -5, 9, -9, 9, 1, 27, -2, -1, -45, 1, -32, 12, 14, 15, -6, -1, 8, 41, 53, 55, 18, 42, 1, 22, 9, -26, -18, -2, -5, 0, 23, -8, -14, 19, -1, -8, -1, -12, -17, -39, 10, -6, -1, 2, 3, 29, 53, 64, 71, 64, 40, 70, 44, 28, 35, 31, 5, 23, 10, -27, -22, 0, -12, -5, 6, -31, -28, -32, 2, -5, -4, 6, 15, 1, 62, 59, 53, 66, 35, 39, 18, 16, 32, 36, 14, 18, 22, 13, -29, -21, -9, -5, 37, -6, 14, 1, 6, 16, -7, 11, -30, 23, 11, 19, -1, -10, 0, -15, 9, 3, 25, 43, 29, 25, 6, 25, 4, 12, -35, -3, 9, 22, -1, 14, -14, 16, 0, 16, -18, 9, 31, 11, 12, 14, -10, 15, 27, 27, 45, 27, 24, 43, 43, 42, 18, 27, -14, -5, -3, 27, -7, -14, 15, 17, 1, 9, 32, 13, 37, 22, 20, 30, 11, -1, 13, 10, -16, 13, 32, 50, 53, 16, 5, -39, -11, -9, -1, 1, 8, -17, -9, -15, -7, 13, 4, -2, 6, -10, -4, -12, -5, -15, -18, -31, 8, 14, 27, 53, 37, 51, 37, 25, -40, -17, -8, 0, 8, 34, 18, -7, 18, 14, 3, -18, -1, -49, -1, -5, 49, 32, 10, 12, 23, 6, 28, 12, 38, 1, 43, 31, 31, -22, 2, -16, 35, 12, 10, -10, -12, -2, -15, -60, -37, -9, 7, 1, -4, 20, 6, -7, 8, -2, 22, -11, 8, -4, 14, 57, 23, 44, -2, 4, 31, 42, -1, -2, 2, -6, -49, -74, -42, -52, -66, -38, 6, -8, 24, 10, -19, 4, 13, -7, 11, -30, -15, 9, -11, 31, 9, 27, 5, 38, -6, -8, 20, -14, -23, -69, -34, 2, -8, -20, -16, -37, -16, 41, 3, 10, 12, 5, -24, -8, -5, -11, -27, -7, -16, -4, -12, -13, 20, -18, 8, 11, 2, -38, -69, -54, -42, -55, -39, -51, -21, -12, -30, -8, -29, -7, -20, -31, -10, 4, -3, 2, 11, 17, 0, -21, -21, -16, 19, 0, -6, -39, -37, -14, -51, -69, -27, -32, -63, -35, -3, -24, 17, -5, -7, -16, -23, -12, -16, -14, -9, -9, -11, 1, -3, 3, -21, 17, 33, 20, -32, -20, -30, -36, -35, 4, -31, -38, -34, -9, -49, -3, 1, 22, 14, -10, -12, -12, 14, 9, 15, 3, -20, 8, 16, 20, 31, 17, -3, -36, -15, -31, -11, -15, 4, -34, 9, 0, -32, -32, -37, 17, -14, -3, 8, -24, 27, 46, 1, -6, 4, 4, 14, -7, 1, -2, -21, 14, -6, -13, -12, 1, 4, -54, -13, -12, -33, -42, -13, -41, -25, -44, -26, 13, 23, 18, 3, -24),
  57 => (18, 9, 13, 2, 16, -14, -18, 15, 4, -13, 16, -9, -14, -5, -14, -17, 9, 11, 2, -11, -19, -4, -8, -3, -3, -12, 2, -7, -8, 8, 6, -17, 7, 9, 18, -20, 14, 9, -6, 13, -16, -4, -18, -26, -13, -12, 44, -4, -13, 1, -23, 5, -14, 17, -17, 14, 16, 8, -7, 11, -2, -14, 4, -19, 17, -17, -16, -35, -1, 29, -8, -17, -7, -34, -53, -74, -17, -3, 10, 19, -14, 4, 2, 1, -7, 15, -7, 3, 7, -18, 5, -13, 5, -28, -45, -4, -18, -7, -19, -21, 7, -26, -1, -8, -14, 3, 18, 33, 4, 6, -5, 7, 18, 8, -18, -13, -19, 13, -8, -22, -14, -2, -39, -14, -9, -5, -7, -17, -23, -9, -4, -2, -7, 12, 7, 19, -21, 0, -6, 20, 10, -16, -6, 13, 0, 20, -28, -2, 0, -19, -15, -5, -27, -12, -25, -10, -30, -22, -12, -12, 30, 21, 34, 38, -21, 12, -11, -9, 15, -8, 8, 4, 2, 10, -17, -13, -42, 26, 12, 6, -16, 8, -32, -38, -11, -19, 11, -25, 18, 3, -9, -21, -30, 12, 1, 6, -15, 4, 13, -13, 12, 5, -1, -10, 2, 0, -15, -58, -38, -9, -35, -9, -9, -21, -20, -23, 4, 2, -19, -15, -23, -3, -8, -7, -2, -10, -12, -16, 18, 17, -10, -10, 1, 2, -14, -25, -28, -21, -17, -15, -20, -28, 2, -14, -2, 11, -24, -53, -34, 2, 20, 5, 2, -9, -5, -15, 0, -3, -46, -18, 2, -17, -6, -23, -45, -45, -61, -27, -26, -17, -27, -15, -18, -10, -2, -47, -35, -26, -26, 20, 17, 0, -4, -12, 18, -4, -66, -69, -62, -28, -16, -49, -25, -32, -55, -22, -37, 3, -10, -44, 1, 4, -42, -53, -17, 16, 28, -17, -1, -19, -4, 11, 19, -10, -59, -59, -41, -33, -40, -48, -30, -6, -20, 11, -5, 25, 19, 9, -4, 7, -22, -26, -18, -7, 12, 23, 16, 5, 0, -9, 10, -2, -15, 9, -5, 0, 6, 6, 23, 14, 36, 31, 11, 50, 13, 25, 6, -21, 19, 28, 5, -7, 38, -4, 2, 19, 3, 15, 31, 12, 21, 42, 43, 56, 45, 73, 41, 45, 37, 31, 41, 34, 31, 16, 22, 33, 19, 11, 29, -11, 12, 15, -16, 10, 4, 9, -14, 9, 28, 55, 54, 48, 41, 28, 47, 21, 13, 41, 31, 54, 33, 20, 26, 24, 25, 39, -36, -34, 17, 22, -20, 11, 19, -21, 17, 15, 46, 40, 33, 40, 27, 30, 17, 32, 7, 23, 40, 27, 13, -12, 35, 21, 5, 27, -21, -51, -11, 9, -20, 20, 1, -3, 37, 21, 26, 24, 17, 49, -11, -1, 7, 33, 17, 4, -2, 9, 6, -4, 11, 11, -15, -2, 1, -43, -10, -5, 12, -6, -15, 16, 11, -12, 17, -11, 7, -19, -53, -68, -50, -57, -44, -5, 12, -21, -40, 2, -10, 8, -16, -15, -31, -15, -20, 12, -2, 5, 3, 10, 22, -30, -35, -70, -54, -47, -101, -119, -61, -49, -51, -30, -19, -48, -30, -31, -39, -26, -17, -31, 9, -8, 35, 3, 11, -15, 12, 9, -14, -3, -57, -46, -56, -62, -40, -57, -55, -44, -39, -11, 7, -18, -24, -36, -12, -25, -29, -29, -7, 4, -35, -20, -12, -4, -20, -8, -23, -14, -52, -68, -8, -3, -46, -42, -28, -30, -20, -28, 0, -62, -34, -13, -36, -35, -28, -13, -3, 6, -19, -33, -19, 6, -5, -5, -13, -41, -19, -59, -14, 17, -25, -48, -60, -52, -35, -23, -6, -47, -59, -19, -47, -40, -31, -26, -22, 17, -12, -48, 18, -3, 15, -14, 2, -42, -59, -70, -8, 33, 4, -10, -18, -16, -43, -25, -37, -11, -21, -13, -29, -64, -21, -38, -26, 3, -7, 8, 13, -8, 19, -6, -22, -13, -24, -9, 28, 60, 60, 7, 0, 17, -10, 13, -5, 28, 34, -32, -37, -47, -29, -43, -45, 2, -19, 5, 8, -10, 10, -14, 18, 32, -13, 6, 36, 91, 52, 11, 44, 26, 60, 42, 35, 5, 30, 3, -10, -2, -39, -23, -15, -8, -37, -36, 3, -9, -10, -9, 13, 38, 36, 23, 17, 20, 18, 18, 27, 13, 29, 46, 12, 8, 16, 21, -4, -21, -7, 8, 23, 5, -19, 12, -17, -10, 15, -3, 17, 7, 16, -3, -14, -31, -28, -18, -8, -21, 17, 9, 25, 12, -1, 24, 9, 11, 18, 17, 42, 49, 41, 5, 0, -8, 6, -10, 10, 17, 8, 12, -28, -55, -47, -14, -6, -16, 16, -1, 7, 9, 28, 53, 60, 49, 47, 47, 52, 18, 56, 37),
  58 => (8, 16, 13, -14, 18, 19, 8, -5, -4, 4, -12, -9, 18, 20, 15, -16, 5, -25, -32, 21, 45, 11, 8, 10, -15, 15, 13, -1, 19, 10, -12, 12, -7, -2, -12, -2, -14, -18, -12, -5, -13, -3, -9, 17, 32, -6, 46, 26, 47, 10, -11, -16, -7, -6, -4, 11, -12, 6, 16, 16, 5, -12, 2, 14, -9, 11, -6, -11, -33, 2, 30, 30, -2, -16, 10, 19, 30, 26, -50, -35, -1, 20, -14, -9, 18, 10, -12, 0, 13, -9, 18, -7, -13, 2, 1, -42, -2, -3, 11, 1, -13, -24, -25, 7, -15, 11, -25, -27, 8, -6, 0, -4, -9, 18, -9, -10, 1, 9, -6, -39, 2, -45, -60, -9, 6, 25, 7, -8, -4, -5, 15, 14, 42, 6, 1, -36, 37, 11, -9, 10, -18, -4, 17, -18, 14, -9, -20, 1, -43, -76, -44, -2, -11, -9, -34, -15, -45, -10, -10, 27, 11, 24, 14, -24, -24, 2, -19, -7, -20, -18, -3, 0, 11, 19, -12, -13, -25, -32, -25, -9, -20, -32, -66, -60, -17, -20, -7, 1, 33, 49, 60, 37, -25, 24, 6, -11, -10, -5, -14, 17, 17, 8, -42, -25, -40, 10, 2, -3, -21, -27, -68, -53, -19, -24, -9, 0, 53, 29, 49, 10, -9, 3, 14, 0, -5, 13, 8, -3, -11, 10, -21, -44, -61, -20, -16, -27, 0, -51, -69, -41, -20, -11, -12, -1, 6, 6, -21, -49, -70, -32, 8, -13, 1, 0, 17, 12, 11, 17, -29, -43, -43, -26, -49, -56, -59, -45, -62, -59, -48, -26, -38, -38, -32, -53, -51, -80, -74, -28, 20, 35, -11, -6, -3, 5, -6, -6, 3, -21, 1, 11, -11, -24, -9, -34, -49, -69, -80, -56, -48, -45, -73, -40, -58, -56, -69, -11, 10, 16, 2, -10, 10, -9, -20, 41, 54, 35, 66, 38, 14, 27, 13, 34, 3, -12, -21, -4, -10, -17, -42, -64, -29, -32, -10, -28, 50, 12, 11, 2, -18, 0, -2, 36, 27, 80, 57, 73, 64, 42, 52, 72, 66, 82, 45, 33, 40, 36, -4, 27, 3, -1, -18, -22, -6, -27, 18, -15, -17, -16, -11, 38, 33, 33, 23, 26, 16, 12, 19, 23, 63, 72, 35, 61, 63, 40, 37, 29, 44, 31, 4, 7, 19, 4, -10, -18, -13, -7, 7, 1, 47, -4, -5, -9, -9, 43, 17, 18, 21, 25, 46, 34, 47, 35, 71, 65, 47, 67, 36, 1, 49, 31, -15, -14, -16, 19, -21, -24, 33, 7, 22, 21, 10, 8, 21, 5, -6, 0, -15, 14, 12, 10, 45, 74, 64, 48, 39, 53, 23, 25, 10, 3, 8, -13, -27, -2, 36, 8, 30, 35, -9, 12, 11, -9, -20, -2, 7, -14, -15, -5, 20, 15, 25, 40, 27, 73, 50, 31, 19, -14, -3, 5, -1, -1, 18, -4, 2, 25, 33, 39, 16, -30, 2, -1, -4, -20, 6, -23, -4, 4, -4, 45, 24, 69, 76, 36, 4, 8, -10, -3, 21, -13, 43, 7, 44, 16, 24, 8, 15, -3, -5, 3, 5, 25, 23, 0, -1, -4, 10, -2, 2, 39, 49, 62, 4, -18, 4, 11, 0, -35, 3, -3, 29, -17, 7, 18, 6, -18, 19, 0, 3, 31, 19, -25, 2, -8, -26, -9, -33, 20, -11, 23, 14, -17, -4, -17, 22, -17, -49, -38, 9, -6, -21, -6, -1, -31, 2, -15, 1, 6, 33, 1, -15, -34, -35, -39, -19, -4, 22, -18, 11, 8, -8, -17, 4, -17, -1, -37, -72, -90, -74, -51, -50, -44, -43, -46, -11, -8, 23, 8, 18, 4, -15, 0, -35, 0, -26, -10, -3, 9, -8, 4, -16, -41, -29, -86, -49, -61, -62, -71, -55, -79, -54, -65, -59, -26, 21, 26, -14, -2, -1, -17, -18, -36, -6, -21, -15, -1, -10, 5, -20, -61, -12, -31, -23, -64, -22, -27, -48, -15, -41, -54, -54, -26, -23, -17, -32, -13, -14, 31, -29, -12, -55, -23, -13, 6, 13, -20, -31, -65, -8, 2, 10, -55, -24, -24, -50, -19, -29, -26, -39, -31, -30, -38, -42, -24, -42, -31, -5, -31, -1, 13, 4, 15, -15, -2, -4, -45, -34, 23, 43, 5, 28, -8, -14, 27, -26, -24, -36, -20, 14, -16, -45, -32, -17, -16, -43, 3, -12, 24, -6, -17, -21, 17, 18, -8, -22, -12, -3, 25, 3, -16, -26, 12, -11, -8, -6, 13, 11, 10, -33, 11, 1, 24, -35, -7, -37, 16, 1, -19, -15, -17, 18, -24, -37, -16, -13, 10, -9, -7, -14, 26, 23, 24, 6, 20, -4, -31, -31, 3, 13, 16, -14, -9, 15, 18),
  59 => (-3, 14, -13, 6, 2, -14, 8, 14, -15, -19, -20, -8, -3, -13, -12, 0, -5, 43, 32, 12, 11, -11, 11, -13, 11, 6, -15, 9, 8, 3, 20, 20, -10, -20, -2, -12, 8, 14, 14, -23, -24, -62, -33, -46, -5, 12, 24, -39, -21, -3, -16, -14, 18, 4, -5, -3, -12, 11, -5, -3, 4, 12, 6, 5, 19, 1, -14, -54, -107, -55, -21, -18, -9, 17, 38, 15, 28, -6, -22, -25, -10, -14, 1, 14, -13, -14, 20, -10, -20, 20, -15, -3, 12, -20, -25, -10, -22, -11, -48, -60, -44, -6, 31, -14, -33, -46, 4, 8, -10, 3, -11, -4, -20, -3, -2, -1, 20, 13, 6, 11, -54, -40, 25, 32, 48, 28, -32, -65, -69, 17, -14, -9, 2, -8, 16, 33, 9, -27, -20, -17, 18, -3, -6, 5, 16, 2, 12, -11, -47, 19, 53, 65, 36, -1, -11, -35, -18, -8, -25, -19, 0, -5, 33, 58, 22, 4, -10, 6, 7, -7, -15, 7, -2, 9, -28, 21, 9, 34, 69, 76, 25, 25, 14, 3, -13, -14, -77, -40, -8, -8, 33, 38, 65, 57, -7, -20, -14, 11, 12, -1, -12, -15, 3, -12, 2, 29, 4, 72, 6, 10, 26, 6, -9, -41, -110, -80, -20, -36, 16, 44, 49, 60, -19, 10, 18, 18, 2, -14, 14, -18, -42, -13, 0, 23, -36, 2, 26, -3, 33, 17, -3, 4, -37, -67, -60, -68, -44, 36, 37, 24, -2, 12, -18, 2, -4, 19, 14, -11, -9, -11, -58, -31, -21, 30, -6, -17, 16, 54, 36, -28, -38, -40, -58, -71, -36, 14, 44, 20, 26, 12, -9, -1, -9, -11, -3, 14, 36, -20, -51, -24, -3, -11, -21, 6, 16, 62, 5, 10, -22, -79, -54, -80, -70, -9, 47, 27, 10, -29, 11, 13, -1, -4, -14, 37, 14, -10, -9, -33, -28, -18, -16, 3, 1, 25, 23, -19, -38, -34, -29, -57, -61, -20, 8, 26, 14, -44, -5, 17, 3, -16, 39, -28, 50, 36, -37, -13, 15, -16, -40, -49, -5, 42, 70, 8, -10, -21, -18, -23, -70, -3, 2, 14, 0, -37, 11, 7, -11, -2, 15, 0, 37, 17, -14, -4, 27, 5, -13, 2, -4, 71, 71, 19, -2, -23, -11, -51, -42, -44, -19, -24, 6, -37, 5, -1, -8, -19, 20, -3, 55, 51, 47, 4, 20, 21, 6, 0, -3, 42, 40, -6, 3, -8, -17, 0, -25, -76, -34, 29, 26, -4, -20, 13, -13, 3, 3, 20, 27, 51, 57, 7, 25, -25, -46, -19, -25, 27, 21, 18, 41, 7, -17, 8, 2, -3, -28, 14, 14, 14, -3, -19, -4, -13, -4, 46, 13, 48, 48, 1, -8, -34, -32, -40, 7, 1, 10, 39, 53, 12, 0, -22, -20, 6, -35, -32, -6, 33, 12, -11, -16, -9, 12, 25, 24, -1, 6, -39, -12, -43, -53, -38, -21, -13, -19, 22, 25, 29, -9, -64, -34, -20, -9, -5, 0, -33, -7, -13, 5, 5, 10, 57, 15, -1, -6, -36, -36, -81, -107, -113, -91, -47, -34, 0, 15, 24, -21, -37, -37, -13, -15, -5, -13, -12, 16, 3, -12, -18, 12, 33, -21, 3, -10, -52, -28, -80, -94, -116, -62, -39, 0, 14, -12, 12, 7, -31, -46, -53, -13, -32, -17, -10, 19, -6, -15, 17, -15, 20, -9, 8, 12, -4, -1, -58, -96, -51, -4, 20, 18, 27, 0, -5, -14, -30, -40, -40, -36, -32, -43, -8, 15, -6, -15, -19, 16, 22, 9, 26, 39, 5, 27, 18, 3, 16, 29, 13, 14, 26, 17, 10, -21, -50, -64, -67, -69, 3, -50, -20, -6, 4, -16, -4, -12, -7, 5, 76, 46, 25, 38, 45, 58, 23, 11, 6, -4, 9, -11, 15, 57, 15, -63, -35, -75, -55, -25, -7, 7, -15, 3, -16, 1, 27, 18, 86, 31, 18, 36, 31, 34, 15, -3, -1, -8, -5, 14, 28, 72, 43, -2, -18, -54, -63, -11, 11, 12, 12, -12, -10, 14, -16, -32, 23, 25, 8, 24, 30, 25, 16, 23, 17, 19, -10, 10, 25, 28, 31, 49, 19, -13, 5, -33, 19, 13, 12, -8, -15, -13, -9, -24, -21, 8, 28, -10, 13, 34, 21, 21, 38, 6, 22, 1, 0, 19, 9, 13, 46, 54, 38, -38, -40, -17, -17, -6, 4, 4, -12, -20, 15, 10, -17, -32, 3, 31, -13, -11, -5, 24, -35, -39, -21, -20, -10, 18, 55, 43, 54, 0, -33, -10, -18, -5, -7, -10, 13, 3, -6, -27, 0, -6, -14, 6, 25, 19, 25, 18, 2, -2, 3, -21, -27, 39, 21, 18, 46, 46, 49),
  60 => (0, -13, 19, -14, -2, -1, 8, 18, 4, -11, 6, 2, -6, 15, 8, -14, -28, -8, -23, -35, -45, -24, -11, 9, 11, -4, 13, -18, 20, -19, 13, 0, -9, -2, 18, -13, 9, 14, 22, -18, 17, 25, 24, -31, 10, -9, 5, -6, -40, -1, 31, 25, -16, -20, 1, -16, -5, -1, 20, -18, 17, -9, -3, -16, 5, -11, 21, 48, 38, 59, 44, 42, 19, 11, 47, 56, 12, 14, -31, -27, 4, -24, 1, -8, -1, -12, 10, -12, -18, -7, -8, -14, 2, 8, -2, 42, 41, 55, 47, 13, -7, 13, -11, -9, 13, -3, -18, 1, -49, -28, -10, 5, 17, 15, -20, -4, -10, 2, 18, -4, -20, -36, 2, 31, 62, 32, 26, -3, 15, -20, -11, 11, -16, -7, 13, -15, -30, -58, 14, 3, 12, 9, 8, 18, 19, 12, -12, -7, -20, -9, 36, 27, 39, 19, 36, 26, 11, -4, 9, 28, 23, 4, -42, -60, -26, -10, 1, -18, -1, -6, -17, -13, -7, 19, -45, 27, 5, 9, 16, 10, 17, 15, -13, -26, -15, 36, 6, 19, 6, -17, -13, -38, 1, -14, 7, -10, 1, -20, -2, -18, 16, -5, 3, 11, 46, 6, -21, -8, 4, -17, -28, -31, 46, 59, 20, -10, 24, 7, 21, 22, 0, 8, 18, 21, -14, -2, 8, 11, 12, 12, 17, 25, 7, -5, -2, -27, -19, -3, -17, 26, 31, 65, 36, 21, 35, 32, 8, 27, 61, 40, 6, 31, 19, -6, 9, -8, -20, 7, 9, 22, 10, -1, 14, 13, 6, 1, 30, 18, 24, 37, 62, 36, 37, 19, 44, 28, 49, 60, 65, 17, 15, 7, -18, 19, 9, 19, 64, 48, 35, 35, 31, 26, 33, 53, 31, 53, 22, 60, 5, -24, 28, 28, 33, 14, 27, 74, 40, 17, -3, 17, -8, -7, -17, 5, 61, 56, 56, 61, 47, 32, 38, 80, 58, 39, 16, 28, 28, 40, 26, 78, 36, 24, 18, 40, 47, 22, -20, -11, 2, 7, 0, -5, 94, 48, 63, 64, 46, 31, 53, 55, 62, 46, 30, 55, 17, 21, 42, 58, 48, -9, -9, 48, 20, 35, -7, -12, 8, -17, 10, 47, 91, 61, 85, 84, 67, 85, 63, 73, 69, 78, 41, 37, 30, 50, 65, 32, 14, -18, -41, 27, 26, 33, -11, -2, 11, 2, -20, 31, 54, 53, 56, 68, 52, 58, 78, 70, 60, 81, 53, 24, 42, 52, 60, 25, 49, 5, -12, 26, 20, -16, 5, 21, -15, 8, -11, 6, -5, 14, 64, 31, 42, 22, 50, 52, 47, 36, 41, 40, 32, 34, 16, 29, 29, 2, -8, 28, 31, 8, -1, 13, 15, 10, 15, 2, 29, 34, 20, 11, 7, -2, 13, 16, 33, 52, 29, 18, 35, 23, 1, 28, -4, 2, 11, -10, 42, 47, 13, -17, 13, 12, 36, 32, 32, 20, 4, 17, -4, -38, -22, 21, 2, 22, -1, 27, -22, 6, 38, 28, 39, 1, 37, 16, 32, 35, -11, -2, 16, 17, 19, 1, 35, 16, -8, -4, -16, -14, -26, 5, 19, 34, 26, 18, -26, 6, 26, 38, 29, 26, 1, -22, 60, 38, -8, 2, -11, 18, 0, 35, 31, -5, -12, 3, -19, 3, -3, 21, 8, -1, 66, 32, 9, 12, 18, 29, 41, 54, 0, -17, 3, 14, -4, -6, -20, -14, -26, 17, 12, -6, -13, -47, -23, 11, 20, 30, 6, 26, 35, 32, 27, 22, 17, 31, 59, 17, 32, -1, -17, -23, 15, -13, 18, 14, -34, 25, 36, -10, -17, -35, 4, 1, -1, 14, 33, 58, 61, 55, 19, -15, 46, 11, 32, 7, 30, 1, -35, -38, -14, -6, -3, -17, 4, 13, 35, 17, -27, -43, 36, 5, 14, -8, 11, 61, 3, 18, 28, 11, 3, 41, 10, 18, 23, 3, -23, -75, 16, 14, -8, -7, -26, 13, 38, -7, -35, 2, -5, 2, -27, -27, 8, 13, 0, 29, 6, 12, 27, -13, 47, 9, 17, 18, 2, -59, 9, 4, 4, 8, 8, -35, 11, 1, 0, -8, 9, -2, -14, 9, 4, 5, -7, 16, 24, 31, 6, 36, 15, 8, 4, 16, 37, -55, 15, -3, 13, -19, -41, -3, 36, -3, -21, -23, 7, 10, -38, -22, -25, -23, -44, 1, -10, -2, 0, 19, 8, 8, 39, 42, 37, -50, 12, 10, -11, -2, -8, 32, 34, -35, -33, -22, -17, -43, -35, -8, -30, 10, 7, 9, 2, -21, -18, -4, -41, -23, 9, 25, -35, -37, -21, 7, 2, 16, -13, 28, 51, 72, 37, 24, 22, 46, 17, 45, 50, 13, 16, 65, 22, 1, -8, -26, -20, -35, -19, -41, -73, -46),
  61 => (9, 14, 5, 8, 2, 17, -10, 5, -20, -1, 12, -19, 11, 4, 1, -16, -24, -12, 19, -9, 19, -10, 7, 17, -13, -18, 14, 10, -6, 11, 9, 0, 18, -13, 1, -6, 7, -11, 5, -8, -4, -11, 11, 10, -3, -14, 16, -35, -21, 7, 6, 9, 8, 5, 0, -17, 8, -4, -20, -12, -20, -14, 20, -2, 6, -6, -28, 6, 1, -20, -41, 18, -20, 5, -6, -6, -24, -82, -60, -48, -20, -20, 4, 11, 7, -18, -1, 10, -5, 17, -8, -17, -5, -24, -31, -28, -61, -76, 15, 8, 12, 10, -8, -13, -27, -82, -63, -32, -47, -18, -15, -8, -19, 15, 11, -9, 9, -6, 20, 3, -1, -35, -66, -64, -78, -29, 14, 31, 18, 5, -7, -29, -27, -28, -33, -15, 3, -12, -10, 3, -16, 8, 10, -3, 15, -12, -6, -8, -34, -61, -86, -67, -53, 3, 21, 27, 37, 14, -18, -26, -29, -37, -22, -39, -7, 12, 10, -2, -5, -6, 16, 20, -1, -3, -20, -20, 12, -77, -52, -76, -32, -4, 15, 5, 20, 19, -38, -26, -37, -4, 14, 6, -13, -8, -9, 3, -6, 9, -14, 14, 11, 16, -20, -54, 4, -43, -44, -50, -22, 1, 25, 39, 23, -11, -36, -18, -12, -17, 9, 18, 1, -54, -9, -10, -4, -14, -1, 3, 11, 14, -32, -28, 12, -26, -45, 18, 20, 57, 55, -13, -28, -32, -39, 23, -2, 8, 41, -4, -7, 26, -8, 3, 18, -19, 17, -3, -20, 2, -14, -20, -38, -29, 15, -5, 28, 38, -22, 4, -10, -10, 12, -4, -4, 0, -4, -5, -20, -9, 18, 10, 3, 10, -5, -6, -16, 10, -54, -25, -31, -8, -18, -5, -16, -11, -7, -24, -26, 15, 4, 0, 4, -17, 21, 3, -43, -41, -3, 6, -18, 5, 9, -19, -3, -15, -70, 15, 22, 13, 25, 25, 28, 6, -14, -32, -15, -2, -19, -8, -4, -17, 23, 23, -15, -7, 12, -8, -10, -21, -19, -17, -7, -8, -37, 47, 29, 25, 48, 45, 7, -3, -29, -36, -40, -25, -16, -13, 6, 1, 13, 23, 21, -34, -8, 6, 1, 9, -16, 16, 17, 19, 4, 41, 11, 4, 12, 0, 22, 1, -14, -36, -36, -1, -34, -23, 29, 19, -10, -14, 11, -5, -41, -3, 0, -8, -17, 17, -22, 20, -10, 12, -6, -18, 1, 5, -28, -23, -17, -44, -19, -7, -10, 20, 27, 13, -3, 23, 34, -18, -53, 22, -2, 6, -11, 14, -38, -45, -41, -29, -54, -44, -22, -55, -31, -43, -21, -49, -1, 37, 50, 42, 20, -16, 12, -23, 1, -19, -40, 7, 7, 15, 12, 12, -42, -82, -62, -28, -81, -68, -37, -35, -27, -14, 46, 47, 59, 44, 17, -6, 13, -16, 17, -20, -35, -5, 4, 25, -5, 8, 15, 2, -18, -113, -24, -47, -66, -28, -25, 0, 14, 28, 66, 49, 28, 63, 25, 14, 33, 18, 4, -20, -48, 12, 60, 54, -14, -14, 9, -13, 7, -64, -24, -31, -3, 18, 66, 46, 43, 57, 19, 19, 48, 59, 15, 20, 14, -27, -67, -55, -28, -16, -3, 12, 13, -2, -12, 3, -21, -10, 7, 20, 38, 58, 83, 63, 61, 37, 22, -8, -9, 11, -14, -45, -70, -17, -74, -48, -65, -47, -30, -26, 9, -17, 20, 6, -24, -2, 41, 60, 64, 55, 65, 53, 25, -1, -5, -34, -17, 5, -54, -68, -61, -36, -76, -28, -5, 1, -20, -69, -20, -14, -13, -8, -11, 38, 21, 41, 77, 60, 22, 17, -8, 5, -15, -3, -37, -46, -61, -76, -48, -34, -13, -25, -19, 0, -1, -38, 15, -20, 8, -9, -18, 6, 38, 26, 39, 46, 19, 3, -8, -27, -36, -88, -77, -118, -73, -34, -75, -55, 1, -18, -13, -21, -15, -16, -15, 10, 8, 6, 39, 41, 0, -21, 14, -24, -27, -40, -52, -80, -71, -123, -118, -109, -94, -64, -70, -68, -18, -34, -13, -11, -8, 0, 15, -6, 7, 7, 51, 45, 35, 6, -48, -57, -81, -68, -76, -107, -79, -62, -93, -102, -78, -35, -33, -32, -18, -35, -9, -19, -21, 5, 2, -9, 13, 7, 1, -4, 25, 14, -48, -82, -71, -52, -38, -45, -32, -42, -25, -80, -46, 14, -19, -28, -24, -17, -20, -29, -2, -12, 3, 10, -15, -1, -5, -7, -39, -21, -1, -55, -46, -65, -22, -31, -31, 5, -20, -59, -14, -14, -28, -10, -48, 15, 14, -28, -13, -8, 17, 16, 0, -6, 4, -23, -11, -19, -16, -37, -16, -32, -48, -20, 5, -7, 3, -24, -20, 19, 4, -6, -1, 19, -14, -12, 22, 3),
  62 => (-8, -10, 20, -5, -10, 19, 19, 7, -9, -8, 3, 16, 15, 2, 13, 27, 48, 33, -15, 17, 31, 1, -1, -4, 14, 8, -11, -17, -14, 8, -7, -10, -3, 11, -12, 9, -11, -1, -32, -14, -8, 15, 44, 36, -10, -67, -20, -11, 26, -1, -20, -1, -9, 3, -1, 20, 10, 7, -4, 10, -8, -16, 18, -3, -10, -38, -45, -31, 25, 20, -2, -53, -31, -38, -31, -13, 38, 8, 8, -14, 16, 12, 0, -17, 17, 5, 2, -19, -11, -14, -21, 8, -4, -74, -13, 4, 6, -19, -66, -42, -91, -58, -44, -14, -8, -35, -2, 12, 37, -9, -10, -19, 18, -18, 17, -6, -8, 14, 18, 9, -68, -20, -13, 2, -50, -46, -25, -27, -51, 0, -25, -12, 1, -32, 5, 17, 67, -12, 7, -20, -18, -18, 20, 10, -20, 4, 15, -69, -19, 2, -14, -62, -43, 2, -7, -12, -9, -16, 28, 32, 29, 27, 35, 24, 11, 17, 1, 4, 12, -3, 0, 7, -3, 18, -12, -71, 26, -3, -43, -24, -34, -31, -25, -21, -9, -16, 1, 8, 26, 51, 29, 34, 9, -16, 12, -10, -9, -6, -10, 6, 17, -8, -24, -5, 1, -1, 25, -14, -16, 4, -2, 2, -10, -31, -2, -16, -1, 23, 39, 16, -8, -21, 33, 24, 0, 5, 4, -15, -19, 7, -26, 15, 0, 64, 21, 14, 10, 9, -11, 24, 10, -4, 0, 15, 6, 16, 61, 21, 19, 31, 41, 41, -13, -5, -8, 17, -10, 20, 36, 55, 33, 69, 29, 31, 17, 5, -19, 8, -8, -31, -19, -12, 3, 11, 15, 1, -10, 29, 20, 45, -20, -20, -13, -16, 1, 61, 73, 68, 52, 56, 64, 20, 16, 4, -16, -11, 17, -20, -6, 2, 5, -27, 8, -36, -17, -18, 43, 35, -15, 8, 15, -3, -1, 63, 116, 4, 40, 41, 27, 28, -29, -15, 3, 6, 11, -3, 12, 14, 13, 29, 16, -15, -2, -23, 12, 50, 5, -1, 1, 1, -47, 35, 24, -19, 19, 32, 29, 37, 48, 32, 32, 15, 15, 39, 6, -6, 30, 29, 10, -23, 0, 5, 36, 21, -6, -19, 17, 19, 11, 18, -17, 3, -8, 27, 54, 103, 80, 41, 45, 16, -2, 48, 54, 42, 38, 20, 23, -1, 10, -14, -14, 38, 0, -9, -6, -6, -28, 10, -10, -28, -40, 1, 5, 50, 53, 67, 22, 31, 65, 7, 22, 11, 5, -8, 36, 19, -17, 15, -23, 41, -10, 10, -18, 20, -8, 10, 27, -23, -75, -55, -43, -23, 25, 0, -15, -23, -17, -1, 23, -18, -20, -1, 2, -18, 10, -10, -4, 16, -13, -16, -15, -9, -33, -40, -77, -65, -124, -93, -127, -127, -88, -57, -73, -64, -50, -39, -17, 4, -32, 1, -6, -16, -7, -21, 16, 8, 13, 6, 18, 12, -28, -44, -120, -103, -149, -146, -106, -135, -123, -115, -97, -77, -42, -41, -28, -6, -9, -15, 14, 1, -25, -3, 10, 29, -17, 0, -17, -4, -30, -45, -58, -46, -30, -50, -23, -36, -35, -58, -32, -10, -24, -35, -28, 18, 27, -4, 20, -25, -9, -19, 4, 23, -9, 16, -10, 4, 1, -17, 13, 18, 46, 57, 25, 16, 10, -11, 0, -1, -17, 20, 31, 40, 33, -12, 18, -9, 34, -4, -35, -12, 12, 9, 16, -5, -50, 2, -15, 22, 31, 48, 22, -1, -2, 9, 0, 3, -28, -12, 10, -26, 13, 16, 6, 28, 8, 24, 11, 5, -1, 9, -15, 4, -35, -31, 10, -25, -4, 31, 17, 23, 50, 37, 40, 27, 30, -4, -16, -16, 0, 6, 8, -33, 9, 4, -9, 31, 10, -14, -13, -6, -34, -41, -15, 33, 10, 25, 7, 36, 42, 18, 11, 13, 10, -24, -12, 2, 14, -35, -39, -44, -7, -22, -2, -30, -7, 17, 0, -4, -17, -69, -13, -28, 13, -27, -3, 13, 14, -59, -48, -11, -39, -32, -25, -8, -65, -43, -55, -27, 17, -25, -44, -24, 7, 1, 19, -1, 17, 9, -44, -14, 4, 10, -25, -36, -24, -22, 8, 18, 2, -42, -32, -23, -15, -32, -49, -33, 48, 19, -24, -45, -8, 13, 12, -19, 16, -10, -11, 18, 19, -22, -46, -30, -24, -20, -7, -12, -14, -55, -8, -36, -24, -28, -61, -65, 31, 27, 2, -49, 19, -13, -10, 14, -11, -15, -13, -34, -13, -57, -46, -27, -40, -26, -14, -23, -6, -59, -30, 17, 21, -3, -75, -89, -21, 41, -35, -23, -12, 1, 14, 13, 6, -13, 12, 2, 3, 1, -9, -7, -6, 1, -10, -43, 17, -37, -31, 26, 51, -11, -20, -3, -24, 10, -3, -40),
  63 => (8, -10, 14, -16, 12, -14, -15, 8, 16, -11, 1, -10, -19, 7, 13, -9, -36, -53, -40, -42, -1, 21, -19, 6, 16, -11, -16, -14, -16, -10, -20, 12, -14, -1, -20, 8, 0, -10, 8, 42, -1, -21, -18, -49, -100, -97, -40, -23, 14, 36, 24, -9, 21, -15, 16, 20, 4, -17, 0, 18, 16, 18, -11, -2, -5, 54, -11, -57, -1, -26, -38, -23, -42, -108, -90, -29, -9, 25, 4, 10, -9, 1, 1, -15, 16, 6, -14, 5, 3, 7, -5, 17, 5, 1, -6, 15, 45, -9, -51, -21, -45, -13, -39, -20, -17, -1, -29, -27, 29, -16, 20, -20, -6, 18, 10, 7, -5, 13, -19, 18, 53, 70, 77, 77, 19, -16, -43, -60, -22, 1, -12, -26, -77, -40, -27, -43, 2, 28, 15, -12, 20, -9, -10, 8, -20, 3, -13, 1, 66, 78, 86, 38, 7, -56, -58, -49, -41, 9, 17, -33, -85, -39, -46, -16, 2, -22, 0, -8, -2, 18, 0, -21, -15, -7, -52, 22, 85, 86, 95, -5, -28, -95, -85, -28, -35, -8, 26, -11, -26, -73, -17, -33, -20, -30, -11, 11, -14, -6, 19, -4, -7, 4, 0, 44, 44, 99, 46, -14, -76, -148, -77, -20, -25, 23, 35, 26, -23, -37, -18, 32, 1, -18, -6, -12, 15, -9, 7, 1, -6, 0, 28, 56, 82, 94, 46, -3, -73, -143, -63, 9, 0, 32, 22, 23, 22, -16, -23, 8, -17, -3, -8, -13, 4, -7, 4, 8, -9, -17, -1, 72, 48, 14, 46, 14, -57, -139, -87, -36, -14, 21, 37, 50, -4, -14, -46, -47, 5, -15, -16, -9, -12, 20, -8, 18, 9, 23, 27, 40, 48, 20, -11, -2, -71, -109, -53, -17, -21, 1, -3, 18, 5, -21, -37, -10, -34, -14, -31, 0, 11, -7, 10, -2, 0, 17, 29, 26, -12, -10, -24, -6, -67, -108, -23, -9, 6, 27, 24, 6, -6, -14, -38, -64, 4, -29, 4, -3, -12, 20, 4, 15, -38, 9, -5, -27, -8, -9, -6, 3, -18, -60, -14, -4, 39, 44, 9, 16, -22, -29, -60, -42, -26, 10, -5, -10, -16, 13, 6, 14, -41, 37, 28, 21, 3, 12, -7, -12, 13, -23, -10, 11, 16, 11, 38, 20, -47, -29, -62, -43, -22, 8, 42, 39, -19, -9, 12, 11, -14, 15, 37, 30, 3, 10, 3, 32, 13, 7, -2, 8, 25, 22, 26, 5, -7, -33, -74, -22, -15, 6, 19, 33, -2, -1, 8, -16, -30, -2, 4, 37, 44, 20, 51, 44, 14, -16, -6, 10, 12, 1, 16, 28, 34, 4, -43, -6, 24, 9, 36, 21, 5, -3, 3, 3, -28, -23, 16, 1, 34, 37, 22, 41, 29, 28, 26, 42, 15, -10, -23, 16, 33, 19, -33, 19, 22, 11, 39, 35, 4, 7, 11, -1, -51, -20, -18, 35, 12, 19, 27, 25, 25, 6, -15, -14, -31, -10, -5, 39, 22, 19, -17, 6, -5, 30, 33, 51, -4, -9, -2, 4, -16, 20, 11, -17, 32, 22, 66, 49, 29, -3, 15, -7, -26, -16, -5, 30, 35, 46, -1, -16, 12, -9, 42, 61, 10, 14, 1, -9, -10, 26, -28, 8, 1, 30, 48, 31, 40, 22, -2, -7, 5, 0, -43, -19, 9, 18, 4, 16, -13, 3, 19, 63, 15, 17, -6, 0, 14, -14, -39, -9, -19, 19, 24, 11, 30, 12, 15, 6, 27, 41, -20, -14, 25, 27, -30, 37, 26, 17, -8, 50, 1, 20, -3, 13, -15, -25, -8, -9, 19, -3, -17, 1, -11, -15, -48, 6, 11, 18, 6, 32, 6, 7, -3, 13, 40, 16, -4, 30, 14, -16, 8, 2, 1, 7, -24, -5, -2, -20, 8, 1, -14, -47, -36, -17, -22, 20, -2, 3, 4, 0, -28, 30, 35, 22, -33, -41, 3, 15, -14, -4, -22, 4, -19, -11, 15, -11, 21, 2, -20, -2, -22, -25, 2, -16, -19, 4, 1, 17, 0, 26, 37, 25, 23, 7, 11, 17, -11, -2, -27, -41, -40, -39, -37, -27, -8, -38, -3, 16, -20, -6, 26, 28, -16, 10, 19, 18, -5, 21, 38, 5, 73, 3, -11, 4, -15, -8, -22, -5, -18, -50, -30, 1, 21, 4, 3, -30, -12, 4, 32, 19, 18, 10, 27, 23, 9, 16, 19, 12, 51, -15, -2, 4, -19, 18, -27, 15, -30, -27, -29, 17, 19, 19, -10, 6, 22, 20, 5, 13, -25, 21, 14, 20, -11, -20, 16, 19, -18, 2, -3, -8, 18, -4, -4, 33, 37, 3, -10, -12, -1, -9, -10, 2, 21, 20, -4, -29, -58, -60, -30, -10, 2, 10, -10, -2, 24, 25),
  64 => (2, 2, -12, -1, -2, -1, 9, -20, -6, 8, 8, 11, -11, 2, -24, -26, -39, -18, 32, 8, 1, 6, -25, -19, 4, -18, -5, -5, -17, 8, 0, -10, -2, 16, -8, 15, 8, 13, -3, 18, 25, -19, -25, -8, 1, -27, 37, -28, 12, -3, -1, -5, -8, 1, 12, -6, 9, 19, 16, -12, 6, 0, 11, 20, -7, -5, 21, -30, -8, -27, -7, -19, 18, 25, 35, 49, 17, 30, 22, -40, -20, -10, 16, -19, -6, 12, 12, -6, -10, -5, 19, 7, 14, -5, 5, 1, 14, 17, 23, 9, 40, 20, 18, 25, 16, 15, 18, -39, 0, 14, -17, 15, 3, -17, -9, -14, -12, 18, 16, 1, 22, 37, 5, 57, 69, 48, 15, -15, 25, 14, -15, -33, 27, 17, 13, -31, 13, -14, 20, 6, -10, -17, 12, -5, -11, 17, 8, -35, 18, -1, -27, 49, 22, 0, 5, -13, 0, 29, -12, -23, -2, -12, -4, -20, 5, 6, 7, -12, -15, -20, 2, 3, 11, 14, 12, -40, -21, -39, -7, -13, 13, 23, 34, -22, 18, -1, -34, 10, -9, 6, -3, -20, 3, -2, 10, 18, -12, 14, 1, 15, 1, 6, -7, -48, -33, -70, -25, -1, 48, -6, 10, 6, -3, -38, -35, -8, -4, -26, -26, 6, 4, -7, -9, 4, -19, -5, 5, -2, -13, -15, -17, -36, -37, -66, -11, 32, 46, 37, 33, 27, -39, -59, -54, -62, -14, -16, -37, -6, -11, 26, 13, 18, -1, 12, 14, 5, -1, -18, 11, -42, -38, -56, -5, 41, 45, 25, 25, 23, -13, -36, -26, -36, 8, -9, 1, -36, -32, 12, 12, -4, -11, 14, -18, 9, 13, 39, -1, -11, -16, -18, 3, 22, 56, 26, 15, 5, -35, -10, -65, -33, -50, -13, -23, -18, -21, -4, -16, -4, 12, 17, 15, 12, -9, -10, -5, -5, 41, 35, 5, 18, 47, 18, 27, 22, -10, -6, -21, -36, -68, -4, -4, -29, -8, 22, -16, -18, -11, 5, -11, -8, 14, 11, -30, -38, 4, 3, 20, 23, 37, 6, -7, 8, 14, -12, -39, -25, -38, -4, -5, -58, -7, 11, 13, 17, 18, -6, -18, 6, 8, 19, -48, -50, -37, -37, -17, 27, 8, 8, -11, -52, -33, -8, -30, -29, -49, -11, 14, -25, -32, -22, -13, -8, 7, 9, 16, -8, -22, -5, -65, -54, -90, -43, 18, -3, 20, 39, -16, -47, -26, -26, -44, -31, -24, -5, 8, -1, -16, -4, -26, -16, 2, -5, -16, -7, -19, 27, -35, -72, -104, -6, -5, 15, 17, 24, -27, -58, -47, -16, 4, -27, -44, -34, 20, 8, -20, -5, -15, 22, -4, -5, -6, -2, 10, 3, -15, -40, -44, -16, -2, 0, -4, 42, -16, -53, -16, -28, -7, -38, -35, -35, 16, 10, -10, -5, -13, 12, 8, -17, 13, 1, 74, -1, 23, 13, -8, -12, 1, -6, 0, -1, -39, -33, -38, -19, -20, -16, -30, -12, -3, -23, -23, -14, 1, 18, 0, 5, 19, 18, 28, 33, 5, 31, 27, -4, 20, 24, 2, -12, -27, -43, -3, -3, 4, -29, -39, 7, 11, -15, -38, -2, -7, 11, 15, 13, 13, -2, 19, 29, 27, 44, -24, 11, 36, 14, 10, 4, 2, -13, -3, 24, -4, -18, -48, -18, 6, -21, -18, -11, 30, -14, -18, 21, 5, 11, -22, -21, 25, 23, 20, 30, 9, -1, 37, 31, -7, -5, 48, 51, 52, 10, 16, 2, -37, -47, -15, -30, 24, -14, 4, -13, -19, 8, -40, 6, 20, 23, -9, 23, -5, 19, 35, -22, 5, -18, 13, 51, 75, 60, 31, 35, -6, -16, -54, -37, 1, 1, 5, 4, 2, -18, 3, -22, -35, 31, 14, 16, -1, 12, 13, -28, -44, -35, -23, 8, 25, 23, 60, 61, 5, 44, 20, 14, 14, 28, 20, -1, 11, 2, 1, 9, -13, -6, 4, -16, -22, 0, -10, -25, -51, -3, -13, 24, -11, -11, -1, 29, 35, 47, 40, 41, 3, 40, -13, -18, -8, -6, 12, -14, -26, -38, -14, 3, 9, 10, -19, -37, -43, -40, 13, -1, -12, -37, -31, 13, 48, -11, 34, 54, 10, 17, -15, -13, 2, -16, 21, -41, -17, -21, -43, 9, 9, 18, -20, -37, -31, -36, -26, 7, -33, -30, -45, -3, 11, -15, 11, 18, 18, 25, 13, 3, -2, -15, -12, 8, -45, -24, -25, -36, 15, 39, 6, -11, -37, -43, 6, 7, 0, -30, -30, -2, 8, 2, -34, 12, 10, -8, 13, -16, 7, 12, -1, 3, -3, -15, -31, -8, 8, 15, -24, -26, -47, -4, -27, -24, -36, -5, 31, -22, -8, 18, -15, 11, -1, 10),
  65 => (14, 16, -1, 15, -11, -1, 5, -6, 2, 19, 6, -16, -19, -3, 17, -18, 7, -34, -22, 10, -29, -58, -4, 14, 12, -9, -20, 2, 14, -18, 2, 10, -4, 10, 19, -12, -11, -19, -16, 15, 1, -17, -14, 11, -10, 11, -24, -35, -38, -25, -20, 11, -12, 18, -10, -14, -17, 0, -7, 9, -3, -8, 13, -12, 1, -10, -12, -9, -4, -30, -42, -32, -34, -30, -54, -60, -71, -67, -15, 16, 16, 17, -9, -14, -4, -9, 19, 3, -2, -5, -6, -10, -3, -5, -34, -51, -51, -40, -47, -18, -35, -40, -36, -20, -1, -22, 14, -2, -22, 18, -20, -4, -11, 19, -16, -12, 18, 0, -17, 20, -2, -16, -16, -26, -35, -73, -58, -45, -18, -6, -19, -1, -29, -4, 32, 30, 19, 11, -9, 15, 4, 3, 18, 10, -18, -10, 15, -7, -17, -60, 2, 5, -13, -4, 0, -3, 2, 2, -2, 11, 35, -2, -2, 13, 8, 9, 17, 17, -12, 2, 20, -2, 13, -14, -13, 13, -3, 27, 60, 29, 42, 49, 41, 14, 39, -2, 20, 62, 42, 19, 35, -12, -4, 21, -16, -5, 0, 20, 8, -19, -11, -16, -1, 7, 40, 32, 3, -20, 21, 54, 34, 42, 38, 31, 28, 25, 33, 50, -9, -6, -36, -34, 2, -2, -18, 2, -3, -8, 3, -3, 32, 20, 12, -17, -14, -52, -40, -40, -8, 5, -28, -7, -11, -3, -25, 12, -15, -50, -14, 3, 9, 25, 8, 16, 21, -20, -4, 7, -6, -2, 2, -15, 6, -5, -31, -45, -23, -49, -80, -82, -18, 4, -15, -10, -84, -79, -47, -5, -4, 15, -20, 9, 5, -8, 15, 36, -20, -27, -3, 48, 89, 88, 48, 28, 54, -14, -56, -64, -36, -40, -24, -15, -50, -60, -47, -21, -14, 15, -14, 10, -16, 6, -14, 24, -26, -14, -29, 25, 51, 49, 42, 30, 44, -3, -30, -16, 6, 35, 30, 14, -19, -4, -30, -22, -20, -11, -17, -1, -4, -3, 30, -12, -34, -29, -5, -27, -35, -15, 1, 3, 13, -54, -80, -26, 20, 33, 17, 4, -13, 0, 1, -16, 3, 17, 1, 2, -14, -14, 4, 25, 21, 24, 23, 6, -43, -28, -16, 4, -3, -51, -27, -3, 30, -8, 42, -5, -25, -30, -3, 4, 0, 37, 9, 8, 20, -17, -16, 6, -5, 17, 16, -4, -46, -55, -65, -11, -32, -14, 26, 16, -5, -17, -15, -14, -31, -36, -29, 2, 1, 36, 8, -2, -10, -3, -38, 5, 5, -43, -28, -32, -40, -83, -98, -79, -70, -28, -12, 33, 5, -18, -12, -19, -31, -66, -69, -42, -1, -48, -16, -8, -19, 4, -44, -24, -85, -53, -57, -25, -52, -61, -71, -50, -46, -13, 3, 22, 29, 40, -4, -5, -36, -26, -9, -13, -15, -16, 14, -18, -16, 8, -35, -32, -40, -18, -22, -12, -11, -26, -25, -47, -21, 0, -15, 3, 35, 32, 3, -4, 6, -1, -14, -14, 8, 18, 16, -5, -18, 2, -22, -62, -53, -32, -55, -26, -22, -10, 0, 10, 18, 2, -6, -7, 25, 36, 38, 1, 35, 7, -1, 18, -3, 3, 14, 10, -7, -12, -3, -14, -54, -107, -87, -70, -22, -16, -14, 19, 32, -12, -44, -34, 3, 23, 37, 27, 23, 11, 38, 10, 52, 36, -12, -15, 1, -19, 4, 1, -38, -92, -85, -33, -31, -30, -7, -16, 51, -25, -14, -22, 18, 22, 20, 17, 29, 52, 54, 42, 45, 61, -21, -12, 12, -15, 48, 45, 9, -8, 25, 6, 31, 12, 29, 29, -7, -3, -12, 28, 30, 11, 1, -16, 22, 67, 32, 33, 61, 51, -2, 11, -19, 5, 56, 53, 40, 40, 37, 25, 30, 24, 22, 16, -6, -5, 11, 47, 46, 50, 17, 2, 42, 32, 27, 9, 34, 67, -21, -5, 9, -17, 73, 59, 50, 46, 45, 24, 24, -2, -6, -16, -12, 0, 40, 25, 11, 54, 31, 27, 39, 13, 9, 16, 4, 24, -4, -6, 15, -19, 35, 46, 16, 1, 1, 8, 26, 30, 33, -4, 21, -10, 4, -23, 12, -4, 12, 21, 23, 56, 28, 15, -2, 19, -20, 11, 12, 11, 19, 47, 53, 26, -44, 0, 29, 7, -17, 18, 26, 52, 41, 30, 41, 1, 3, -6, 8, 27, 25, 15, 11, 34, -5, -10, 3, -17, 7, 6, 32, 34, -22, -21, -27, 11, 6, 38, 64, 51, 51, 48, 27, 21, 14, 16, 34, 16, 15, 1, 41, 31, 12, 11, -7, -2, -19, 2, 2, 36, -24, -4, -6, 19, 29, 36, 23, 0, 17, 29, 20, 16, 10, 32, 38, 35, 4, 12, 19, 60),
  66 => (-4, 11, 19, 15, 8, 3, -20, -4, 4, 3, 7, -4, 5, -4, 39, 57, -3, -24, 5, -4, -18, -8, 3, 11, -15, 14, -10, 13, -18, -15, -9, -16, 8, -10, 6, 3, 6, 16, -5, -24, 17, 56, 67, 77, 68, 37, 49, 32, 19, -7, 14, 10, -7, 8, 4, 19, 8, -3, -12, 5, 2, -2, -8, 7, 4, 12, 4, 51, 28, 30, 1, -19, -39, -11, 8, 36, 31, 36, 17, -23, -9, -8, 12, -11, 4, -10, -6, 19, 15, 4, 11, 6, 16, 30, 37, -33, 4, -38, -2, 13, 2, -26, 7, 6, 9, 13, 2, 2, -19, 5, 5, -2, 11, -3, -4, 5, -12, -13, -19, 15, 24, -2, 10, 47, 2, -23, -6, -3, 16, 8, 29, 14, 19, 5, -1, -26, 5, -4, -5, 14, -6, -18, -10, 14, -12, 5, -19, -7, -32, -31, 27, 45, 4, -9, -25, -14, 13, 26, 21, 13, -4, -3, 5, -4, -26, 19, -14, -9, 3, -12, -1, 16, -3, 11, 15, 29, 33, 20, 3, 8, -9, 4, 18, 9, 16, -9, 19, 31, -13, -28, 24, -31, -31, -32, -4, -13, 13, 3, 21, -14, -13, 14, 4, 24, 39, 52, -6, 23, 17, 17, 38, -5, 7, -2, -9, 11, 13, 2, 3, 9, -64, -32, 3, -13, -5, -4, -20, -7, -8, -11, 30, 51, 48, 59, 32, 21, 43, -6, 5, 15, -24, -15, -23, -7, -18, -33, -26, -58, -72, -21, 7, 8, -15, -4, 7, -2, 18, -4, 16, 11, 24, 27, -7, 39, 50, 33, 37, 2, -1, -25, -29, 8, -8, -14, -20, -73, -86, -33, -36, -12, 9, 11, 3, -19, 0, -36, -28, -60, -49, -21, -4, 10, 19, 15, 52, 12, -2, -35, -26, 13, -20, -19, -16, -60, -106, -44, 27, 58, 15, 0, -12, -16, 14, -44, -83, -139, -107, -25, 37, 35, 1, 39, 50, 20, -1, -9, -6, -23, -24, -32, -8, -20, -19, -28, -12, 70, 13, -18, -1, 5, 24, -22, -89, -109, -95, -32, -28, 16, 13, -9, 9, 20, 43, 18, 25, 3, -5, -32, -13, -24, 4, -16, -41, 11, 16, 18, 14, -6, 4, -32, -68, -122, -136, -78, -22, -14, 9, 27, 7, 43, 59, 20, 35, 1, -28, 6, 17, -11, 8, -14, -13, 11, -18, 0, -10, -14, -3, -19, -53, -72, -105, -119, -72, -26, -29, 0, 1, 22, 58, 62, 35, 12, -19, -27, 16, -15, -13, 14, -9, 43, -11, 6, -8, -2, -17, -28, -71, -106, -91, -71, -91, -90, -59, -26, 3, 33, 63, 44, 15, 14, 8, -12, -28, -21, -14, 24, 19, -4, 10, 15, -2, -11, 3, -35, -62, -58, -67, -27, -70, -114, -129, -27, 1, 30, 34, 22, 54, 38, 18, 6, -22, -9, -2, -3, -15, -15, -6, -10, 6, -6, 8, -37, -27, -11, -44, -79, -73, -109, -124, -78, -12, -19, 18, -1, 32, 10, 19, 17, 26, 29, 10, -1, -8, 21, -6, -18, -19, 19, -29, -5, -32, -38, -29, -47, -59, -117, -179, -48, 7, -31, -9, -3, 20, 40, 27, 37, 17, 35, -5, -34, 6, -25, 1, 11, -8, 16, 1, -14, -30, -23, -48, -52, -86, -80, -139, -31, -5, -54, -12, 7, 8, 24, 5, 80, 13, 38, -5, -6, -5, 4, -14, 4, 0, 5, -16, -10, -13, -26, -38, -41, -45, -81, -127, -49, -12, -51, -52, -3, -12, -17, 23, 75, 40, 22, 32, -8, 40, 34, -10, 6, -11, -16, 9, -14, -43, -32, -15, -38, -29, -91, -111, -40, -46, -41, -21, 2, -19, -11, 3, 39, -8, 8, 3, -7, 20, -37, 10, -19, -3, 7, 9, -16, -14, -38, -36, -32, -46, -61, -103, -105, -70, -42, 4, -8, 17, -41, -25, 14, -22, 25, 2, 10, 9, -48, 14, 15, -11, 12, 5, -20, -7, 7, -15, -5, -43, -3, -50, -74, -93, -33, 12, 10, -22, -24, -6, 4, -20, -1, 27, -9, 26, -19, -18, -1, -17, -8, 20, 16, 19, -11, -10, -23, -17, -34, -66, -71, -80, -53, -29, 3, -16, -40, -1, -21, -36, -10, 36, 14, 24, -32, 6, -1, 19, -20, 16, -14, -19, -14, 3, -18, -3, -23, -19, -84, -71, -44, -13, -33, -25, -16, -13, -24, -30, -27, -17, 16, -20, -29, 5, 7, -20, -5, 19, -3, 2, -4, 13, 2, -33, -36, -40, -15, -30, -8, -1, 9, -2, -30, -28, -25, -36, -19, 36, -1, -40, -29, 17, -8, 1, -12, 2, 3, -4, 11, 1, 18, 2, -6, 1, 4, -35, 21, 70, 19, 5, -25, 2, -3, 3, -13, 27, 42, 1, -9),
  67 => (6, -13, -15, -6, 5, -11, -12, -19, -20, -4, -10, 3, 11, -5, -29, -61, -49, -64, -43, -78, -39, -29, -5, 16, -19, 18, -6, 12, 14, -10, 6, 0, -7, 11, 2, 20, -14, 13, 27, 65, 56, 14, 12, -20, -8, 9, 0, 1, -11, -16, 11, 22, 12, 5, -21, 10, 18, 8, 6, 16, 4, -13, -14, -15, 3, 75, 42, 53, 68, 57, 38, 49, -9, -7, 10, 39, 7, -16, 5, 41, -8, 30, -5, 10, -6, 8, -16, -5, 18, -17, 17, 4, 54, 17, 42, 57, 84, 45, 24, 24, 10, 5, 11, 43, 36, -14, -28, 13, 6, 3, 11, -9, -15, 5, -10, -3, -20, -17, 3, 48, 29, -16, 35, 36, 41, 34, 44, 13, 17, 26, 26, -20, -6, -11, -28, -35, -28, -35, -7, 2, -15, -12, 1, -6, 7, 13, 16, 63, 55, 12, 4, 32, 36, 59, 41, 14, 10, -13, 21, 18, -26, -39, -36, -5, -22, -55, -17, 8, -20, 12, 7, 10, 4, 13, 43, 72, 21, 16, 18, 48, 42, 35, 12, -4, 6, -14, -35, 21, 13, 13, 49, -3, 7, 31, 13, 9, 3, -3, 7, -9, 18, 2, 73, 44, 35, -11, 22, 27, 27, 18, 28, 4, -26, -12, -53, 0, 14, 15, 35, 1, 30, 50, -6, -1, 19, 13, -6, -9, 20, -5, 20, 3, -1, -3, 54, 58, 56, 44, 23, 12, 4, 38, 1, 32, 52, 8, -4, 44, 65, 22, -25, 19, -1, 19, -14, 0, -2, 19, 10, -9, -25, -18, -8, 17, 38, -3, -5, 3, 16, 16, -8, 29, 79, 70, 51, 71, 63, 62, 43, -1, -15, -18, 13, 0, 5, -22, 5, -8, -40, -43, -56, -32, -4, -33, 3, 10, 23, 16, -2, 10, 58, 68, 38, 36, 10, 10, 28, -38, -2, 3, -6, 20, 0, -17, -13, -31, -69, -56, -47, -14, -4, -10, -6, -2, 10, -9, -12, 13, 14, 22, 51, 46, 4, 19, 26, 1, 17, 10, -17, 6, 35, 41, 26, -44, -18, -3, -12, 31, 24, 21, -19, -3, -18, -11, -18, 8, -14, -7, 19, 27, 20, 35, 57, -35, -13, 13, -5, 3, 64, 46, 58, -11, -9, 23, 3, 47, 20, 27, 8, 25, 5, 31, -10, 8, 9, 3, 11, 39, 1, 36, 33, -7, -18, -11, -7, 9, 19, 33, 66, 17, 27, 19, 13, 44, 24, 34, 58, 32, 23, 64, 33, 31, 29, 34, -29, 24, 46, 29, 21, 3, -13, 14, -5, 12, 7, 63, 17, 30, 25, 42, 36, 20, 38, 24, 35, 29, 36, 63, 43, 43, 71, 63, 16, 16, 17, 47, 8, 7, -19, 10, 4, 8, -1, 67, 22, 32, 56, 38, 77, 30, 24, 24, 48, 42, 51, 50, 63, 69, 65, 109, 26, 14, 30, 26, -10, 46, -19, 10, 3, 18, 6, 24, 77, 49, 55, 19, 48, 47, 35, 37, 58, 50, 85, 81, 66, 44, 47, 57, -2, 12, 59, 72, 21, 25, -21, -12, 10, 15, 16, 9, 42, 57, 39, 43, 48, 67, 63, 68, 34, 51, 69, 18, 57, 40, 21, 28, -7, 9, 21, 31, 15, 48, -5, 0, 11, -9, 16, 17, 32, 28, 59, 54, 63, 39, 55, 78, 70, 42, 53, 78, 51, 14, 0, 38, -5, 25, -12, 24, 11, 44, 1, -5, 20, -20, 21, 41, 72, 50, 59, 53, 36, 71, 59, 35, 61, 38, 52, 53, 33, 17, 13, 19, 29, 8, 10, 41, -19, 50, 13, -2, 4, -4, 10, 82, 76, 55, 75, 37, 26, 24, 34, 26, 36, 36, 33, 37, 53, 40, 0, 26, 3, -3, 32, 26, 17, 22, 15, 3, 9, -4, 62, 41, 52, 35, 50, 14, 26, 33, -18, -35, 20, 24, 22, 33, 15, -16, 7, 17, -20, -18, 27, 49, 20, 17, 12, -21, -16, -13, 15, 27, 56, 14, 8, -12, 14, -18, -38, -13, -4, 40, 39, 6, -5, -4, 41, 3, -17, -15, 6, -4, 22, 17, -11, 18, -19, 20, 6, -8, 1, 18, -19, -23, 10, -14, -11, -8, 5, 18, 0, 33, -14, -17, 9, 21, 23, -24, 1, 12, 47, 41, -9, 1, -3, 12, -44, -8, 2, -7, -4, -25, -14, -8, -38, -25, 7, 13, 13, 2, -42, -37, 3, 39, 8, 35, 12, 22, 25, 5, 17, 6, 6, 5, -33, 39, -23, 1, -11, 7, -40, -73, -49, -7, -7, -15, 17, -5, -7, -27, 23, 36, 3, 9, 3, 9, 24, 24, 0, 6, 9, 15, 1, 46, 41, 37, 50, 8, 32, 11, 35, 28, 12, 24, 21, 13, 25, 3, 3, 9, 17, 3, -13, 26, -23, -6),
  68 => (4, 2, 7, 9, -3, 5, 12, 12, 17, -8, 20, 0, 18, -10, -12, -15, 5, 12, -17, -18, -5, -17, -13, 12, 3, -4, 15, -1, 9, -8, 0, 16, -18, -3, -14, 20, -1, 3, -2, 6, 17, 29, 37, -8, -10, 18, -17, 3, -23, 2, -5, 1, -15, -19, -20, -1, 0, 20, 14, 13, -7, 17, 11, 14, 7, -1, 5, 4, 17, 29, 25, 23, 25, 8, 19, -14, -38, -17, 12, -10, 7, 12, -9, -19, -6, 11, -14, 16, -1, -9, -11, 17, 14, -10, 7, 45, 5, 20, 28, 9, 17, -9, -5, -17, -35, -33, -37, 1, 4, -9, 10, 12, -15, -1, -4, -19, 18, -17, 7, 17, -24, 1, 23, 35, -2, -34, -14, 38, 15, 6, -9, -39, -25, -51, -35, -38, -35, 2, -12, 11, 15, -15, 2, 7, 1, -7, -7, -7, -3, 6, -17, -22, -36, -1, -8, 24, 29, 8, -26, -11, 2, -20, -41, -10, -28, 10, -15, 16, 12, 10, 10, 9, 1, -13, -12, -14, -9, -8, -17, -13, -22, 13, 19, 10, 20, 21, -16, -7, -34, -9, -43, -34, -21, 23, -10, 10, -8, -12, -12, -10, -4, 13, -19, -24, 22, 25, -13, -4, -12, 8, 31, 22, -11, -49, -44, -11, -15, 3, -11, -68, -23, 14, -5, 6, 17, -11, -4, 5, 8, 8, -42, -23, 7, 5, 2, -21, 6, 8, -6, -17, -23, -47, -34, -17, -26, -2, -5, -18, -4, 20, -20, 15, 18, -18, -18, 6, -15, 13, -17, 23, -7, -22, -16, -38, -14, -7, 6, 0, -36, -20, -39, -28, -22, -15, -27, -14, 40, 35, 0, -14, -7, 2, -19, 1, -20, 8, 5, -37, -21, -13, -5, -30, -19, -13, -26, -29, -19, -30, -9, -24, -32, -35, 0, -7, 9, -3, 9, -9, 8, 20, -2, 2, -19, 3, -7, -41, -30, -28, -28, -56, -35, -29, -11, -56, -42, -51, -50, -20, -9, -18, -13, -14, -6, 38, -8, 2, -2, -15, -13, 21, 5, 2, -53, -42, -43, -60, -11, -45, -40, -38, -53, -16, -31, -40, -26, -17, -4, -39, -26, -7, 15, -4, -58, -6, -17, 0, -17, -12, 10, -41, -48, -56, -64, -55, -30, -38, -13, -34, -59, -46, -32, -31, -42, 7, -4, -53, -39, -31, -2, -15, -57, -31, 11, -20, -17, -7, -18, -16, -42, -28, -55, -93, -42, -48, -41, -32, -30, -53, -62, -7, -20, -27, -24, -22, -16, -20, -3, -26, -9, -13, -16, -12, 16, -21, 7, 7, -19, -23, -51, -48, -38, -61, -36, -44, -50, -45, -56, -5, -17, -9, -3, 10, -2, 10, 3, 32, 3, 52, 12, -8, 18, 15, -14, 16, -2, 1, 26, 12, 0, -27, 4, -14, -15, -16, -15, -5, 9, 35, 39, 2, 19, 25, 36, 36, 24, 57, 6, 12, 12, 4, 27, 42, 7, 63, 39, 41, 50, 61, 88, 69, 76, 27, 42, 61, 42, 34, 19, 24, 20, 24, 26, 32, 22, 49, 7, -9, 15, 6, 44, 47, 54, 60, 62, 52, 69, 66, 84, 58, 54, 68, 54, 44, 23, 37, 32, 12, 22, 30, 33, 17, -11, 63, 2, -18, -19, -6, 69, 45, 50, 46, 36, 67, 42, 28, 38, 56, 25, 69, 49, 60, 31, 2, 43, 3, 9, 36, 18, -7, 15, 76, 16, 13, -6, -6, 57, 28, 69, 29, 37, 49, 24, 27, 44, 49, 36, 64, 43, 26, 5, 7, -3, 22, 38, 36, 1, 2, 7, 42, -1, -7, 4, 15, 47, 2, 23, 28, 20, 8, 14, 39, 74, 44, 36, 64, 40, 29, -1, 16, -12, 5, 25, 7, 33, -4, 41, 89, -9, 3, -7, -17, 69, 31, 7, 10, 28, 36, 24, 40, 59, 24, 40, 22, 23, 57, 21, 30, 39, 38, 0, 41, 11, -11, 47, 55, -13, 19, 5, -9, 67, 40, -2, 8, -3, -11, 0, -15, 14, 24, 27, 5, 36, 47, 35, 36, 35, 32, 31, 59, 29, 4, 68, 59, -12, 13, -11, -12, 5, -12, -9, -32, -29, -35, -22, 19, -9, -5, 4, 0, 11, 2, 34, 16, 18, 52, 32, 20, -4, -26, -13, 37, -13, -4, -13, -6, -18, -29, 24, -18, -24, -41, -15, 5, -16, -25, -5, 5, -5, -28, 8, -17, 37, 40, 26, 9, 9, -27, 12, -9, 11, 0, -5, 8, 9, -19, -1, 9, -36, -36, -9, -28, 6, -37, 2, -16, -31, 1, -4, -24, 36, 58, 24, 28, 50, 9, -17, -3, -3, -8, 15, 13, 1, -41, -12, -20, -26, -3, -32, -13, -13, 12, -22, -33, -35, 5, 17, -1, 10, 7, 27, -1, 15, -8, 15, -4),
  69 => (4, 14, 17, 7, -18, -10, 20, 15, 4, 5, 21, -10, 6, -1, 6, -24, -29, 24, -28, -27, 17, -4, 4, -8, 7, 19, 4, 5, 13, -18, 13, 14, -3, 3, -11, -7, -4, 14, 17, 3, 44, 7, 19, -16, -44, -30, -50, -35, 52, -12, 5, -9, 1, -15, 12, -20, 7, 9, 10, -9, 12, -13, -9, 2, 13, 35, 30, 27, 71, 24, 24, -17, -44, -82, -59, -51, -32, -81, -26, 6, 4, 1, 19, -6, -11, 17, -1, -12, 7, 6, 1, -4, 22, 31, -7, 6, 18, 44, 10, 27, -8, -27, -35, -32, -63, -75, -54, -10, 22, 21, 19, 1, 20, 10, -8, 0, -6, -1, -13, 13, 43, -63, -27, 15, 29, 19, 41, -2, 16, 23, -28, -47, -69, -61, -30, -37, 25, -18, 9, -13, 20, 17, -13, -13, -19, 20, 30, 57, -20, -18, 14, 49, -2, 16, -14, 32, 32, 47, 2, -27, -30, -72, -51, -12, 16, 45, -11, 2, 4, -3, -1, 7, 6, 0, 40, 40, 41, 27, 48, 43, 21, 3, -23, 7, 36, 63, 45, 22, -1, -96, -50, -15, 22, 37, 17, -16, 7, 5, -3, 8, -19, -19, 79, 33, 121, 75, 59, 40, 20, 13, 6, 12, 22, 10, 3, 9, 12, -67, -72, 20, 44, 17, -20, -11, -2, -12, -18, 10, 12, 9, 69, 33, 110, 63, 44, 63, 40, 19, -40, -39, -1, 8, -7, -48, -20, -79, -91, -19, 40, 34, -13, 9, -13, -18, 10, 17, -21, -10, 27, 9, 48, 61, 37, 52, 70, 6, -48, -2, 17, 31, -7, -46, -37, -49, -82, -43, 12, 5, -22, 22, -13, 14, -12, -13, -15, -15, -31, -8, -31, -15, 38, 28, 38, -32, -75, -58, 0, 27, 24, -28, -41, -51, -79, -34, 13, 25, -17, -16, 6, -7, -5, -6, 20, -37, -50, -40, -56, -2, 1, -7, 17, 9, -45, -59, -36, -2, 31, 15, -21, -47, -66, -74, 30, 5, -15, -11, 11, -11, -9, -19, 22, -66, 11, -39, -64, -37, -37, -31, 11, 15, -37, -19, -10, -29, 27, -8, -29, -59, -91, -67, -6, 5, -18, 22, 14, -15, 16, -14, 35, -28, -19, -75, -78, -72, -67, -25, 0, -26, -35, -19, 38, -7, 23, 16, -21, -52, -77, -60, -13, 10, 6, 52, 9, 17, 10, -7, 19, -30, -54, -64, -46, -73, -77, -38, -33, -32, -12, 4, 19, 10, 11, 10, 40, -4, -35, -16, 7, 6, 9, 38, 15, -3, 10, 16, -12, 0, -20, -46, -12, -37, -41, -42, -48, -37, -19, -6, -10, 42, 20, 25, 27, 83, -9, -43, -2, -9, 9, 30, -5, -1, 19, -9, -12, 27, -12, 29, 31, 7, -33, 12, 4, -24, -2, -9, 8, 36, 37, 13, 44, 68, 34, -19, -6, -14, 39, 53, 12, -14, -2, -20, 13, 5, 10, 24, 46, 62, 4, 30, 9, -9, -18, -5, 15, -2, 2, 26, 44, 57, 20, -46, -40, -16, 44, 63, 3, 7, 13, 12, 43, 52, 14, 21, 42, 29, -8, 5, -5, -6, -1, 22, 6, -3, 26, 43, 50, 70, -4, -36, -39, -28, 3, 29, 5, 18, 15, 19, 44, 29, -10, -25, 16, 24, 2, 17, 6, -5, -3, -10, 11, 5, 4, 16, 47, 18, -1, -24, -39, -39, -8, 24, 8, -5, -11, 17, 82, -14, -48, 5, 2, -2, -32, 8, 8, 24, 6, 0, 12, 33, 31, 28, 41, 27, 12, -58, -48, -1, -41, -20, -6, 14, -1, -6, 32, 18, -29, 25, 4, 26, -12, 9, 1, 28, 20, -36, -4, -16, 26, 43, 5, 30, -2, -20, -52, -6, -40, 2, -18, -14, 10, 6, 55, -33, -39, 7, 20, -24, 12, -24, -5, -29, -19, -21, -35, -48, -56, 24, 37, 35, 3, -30, -56, -20, 10, 33, 10, -19, -4, -10, 2, -23, 0, 30, -17, 12, -15, -57, -40, -51, -61, 7, -17, -16, 22, 10, 40, 56, -9, -47, -55, -24, 20, 74, -3, 6, -16, 20, 8, 19, -10, -15, -45, -7, 6, -19, 9, -34, -25, -40, -32, -7, 51, 36, 45, 75, 11, -45, -72, -39, 22, 31, -14, 18, -2, -15, -13, 38, 30, -8, -45, 3, -15, 0, 3, -10, -19, -41, -68, -3, 25, 8, 5, 23, 5, -23, -46, -53, 15, 39, 15, -5, -20, -16, -6, 61, 54, 26, -35, -29, -22, -7, 3, 3, 19, -6, -46, -70, -44, -2, -15, 4, 2, -2, -11, -4, 15, 24, 5, 2, 18, 1, -2, 25, 63, 47, 23, 30, 10, 12, -2, 0, -12, -8, -37, -26, -9, 3, -18, 10, 79, 56, 35, -1, 19, 27),
  70 => (-14, -1, 16, -18, -17, 13, 5, -1, -5, -7, -1, -19, 0, 2, -30, 14, -5, -30, -24, -24, -9, 12, 13, -18, -19, 7, 14, 20, 8, 11, -3, -4, 4, 3, 9, 4, 14, 20, -17, 8, 20, -1, -17, 37, -16, -18, -10, -12, -2, 3, 16, 4, 35, -2, 6, 8, 12, -3, 19, 12, 11, 14, 18, -6, -15, -13, 11, -1, -23, -19, 5, 5, 2, -9, -3, -21, -19, 10, 38, 20, 37, 3, 5, -5, 7, 7, -18, 14, -9, -15, -20, 5, -2, 17, -27, -36, -34, 0, 18, 18, 10, -7, 5, -42, -32, -5, -17, -21, 2, 10, -11, -13, -13, -3, -2, -20, 0, -14, -7, 6, 19, 17, -2, 27, -3, -42, -25, 15, 35, 28, 13, -15, -7, -11, -5, -31, -29, -9, -17, 14, -12, 18, 20, -18, 11, 19, 9, 12, 12, -11, 43, 36, -16, -7, -9, 41, 23, 15, 1, -11, -39, -47, -22, -32, -52, -23, 3, 9, -18, -14, -19, 13, 0, -20, -19, 34, 22, 16, 51, 42, 11, 1, 44, -4, -34, -20, -24, -39, -31, -37, -39, -23, -14, -28, 7, -7, 20, -5, -12, -3, 15, -7, 9, -31, 19, 41, 40, 69, 32, 30, -20, -39, -23, -41, -3, 7, -35, 0, -27, 15, 23, 10, -7, -3, -17, -2, -11, -15, 0, 18, -9, -4, 42, 29, 41, 55, 6, -34, -12, -25, -14, -44, 31, 4, -9, 20, -2, 25, 65, 15, -16, 2, 3, 5, 19, 1, 11, 2, -46, 21, 65, 24, 35, 11, -34, -57, -32, -26, -1, -4, 30, 34, 21, 10, 12, 35, 29, 19, -15, -3, -11, -19, 1, -3, -15, -17, -49, 45, 42, 48, 14, -40, -75, -78, -22, -27, -30, -15, -5, 18, -10, 11, 9, 23, 40, -3, -20, -16, -9, -5, 14, 8, 2, -69, -27, 49, 4, 3, -24, -29, -65, -73, -16, 6, -31, 11, -2, 15, 23, 28, 16, 18, 37, 8, -21, 7, 8, 3, 10, -18, -14, 0, 15, 14, -32, -57, -26, -3, -48, -65, -1, -32, -31, 10, -17, 4, 26, 3, -4, 37, -12, 1, 2, 2, -8, 20, -5, -1, 4, -34, -2, -38, -57, -16, -26, -1, -59, -19, 20, 1, 31, 17, 22, 12, 33, 10, 25, 31, -20, -19, 4, -12, -3, -9, 12, -13, -35, -38, -14, -26, -64, 4, -22, -24, -8, 18, 40, 11, 50, 31, 49, 25, 34, 20, 47, -8, -33, -20, -44, -15, 5, 18, 12, -11, -33, 4, 42, -10, -17, -2, 36, 50, 45, 47, 25, 6, 36, 33, 22, -8, 40, 26, 38, 20, -22, -35, -31, -41, 17, 14, 4, 19, -10, 10, 30, 43, 14, 34, 31, 10, 29, 25, 28, 23, 44, 26, -17, -8, -8, -25, -8, -13, -48, -35, -17, 4, 6, 0, 14, 15, -15, 26, 24, 41, 27, 33, 39, 17, 31, 35, 42, 11, -4, -30, -47, -27, -52, -62, -48, -21, -48, -42, -26, 21, -2, -7, -12, -8, 12, 24, 9, 38, 59, 15, -3, -13, 13, -14, 8, 2, -25, -17, -25, -45, -46, -36, -58, -51, -44, -44, -5, -15, -9, 4, 1, 8, 25, -4, 0, 23, 2, 3, 25, 6, -24, -55, 3, -22, -15, -4, 6, -50, -19, -50, -46, -41, -32, -52, -41, 13, 20, 10, -10, 3, 20, 19, 8, -25, 8, 9, 19, -45, -70, -37, -51, -50, -59, -21, -2, -37, -2, -28, -32, -42, 2, -23, -40, -27, -3, -18, 6, -10, 23, 42, -6, -6, -10, -10, -21, -33, -84, -76, -68, -50, -28, -29, -24, -32, -24, -29, -33, -32, -30, -18, -25, 7, -18, -2, -3, 7, 29, 20, 1, -3, -54, -57, -22, -23, -75, -81, -72, -32, -24, -32, -12, -35, -25, -20, -45, -6, 1, -25, -33, -4, -1, -16, -7, 16, 17, 48, 27, -17, -31, -23, 4, -13, -15, -53, -36, -30, 2, -62, -31, -37, -46, -17, 9, 3, 6, -4, -46, -6, 12, -13, 1, 21, 29, 24, 27, 34, -19, -27, -5, -24, -33, -21, -13, -29, -7, -21, -53, -7, -15, -23, -3, -20, 7, 20, 18, -2, -6, -13, -6, 5, 1, -7, -6, -15, -19, 4, -3, -26, -13, 4, -1, 38, -29, -13, -15, -21, -29, 3, 23, -3, 3, -1, 3, 0, -13, 10, -20, -9, 14, 6, -15, 2, -13, -8, -14, -4, -16, 13, 3, -25, -14, -5, 21, -1, -5, -4, 28, 1, 15, -2, -16, -1, -11, 11, -18, -17, -13, -2, -20, -6, -1, 19, -7, -19, -16, 2, -7, 20, -15, -7, 5, 20, -12, -2, -12, 7, 1, 7, 11, -8),
  71 => (-7, -15, 0, -12, -14, 12, 15, 18, -18, -14, -11, -9, 9, -1, 11, -26, -21, -72, -49, -40, -21, -36, -46, -19, 15, 4, 2, -11, 10, 18, -6, -9, 7, 14, -19, -10, 14, 11, 40, 71, 48, 30, 40, 10, 34, 19, 8, -21, 27, 8, 14, 23, -3, 20, 14, -15, 5, 6, -17, -16, -15, -17, -5, -8, 7, 54, 23, 91, 56, 13, 6, -19, -45, -15, -11, -24, -18, 19, 7, 44, -7, 2, 18, 4, 16, 14, -8, -10, -14, -12, -7, 17, 81, 44, 71, 62, 24, -4, -9, -32, -62, -30, -35, -10, -27, 44, 41, 26, -29, 13, -7, 9, -2, 17, 0, -17, 5, -19, -13, 43, 56, 29, 29, 44, 34, 2, -21, -60, -16, -1, -13, -10, -22, 0, 15, 17, -47, 3, 7, -16, 19, -20, 20, 10, 9, 1, 30, 28, -11, 8, 32, 38, 26, -8, -2, -29, -18, 0, 9, -4, 10, 13, 16, 21, 7, -14, 10, 15, -10, -18, 14, -1, 13, 13, 25, 45, 15, 38, 32, 6, 24, 48, 9, 9, -9, 1, 13, 7, -3, 9, 38, -20, -8, 16, -19, -1, -19, 9, 4, -1, 6, 5, 44, 82, 36, 3, -26, -12, 38, 36, 31, 12, 30, 25, 7, -23, -2, -5, 9, -7, -22, 11, 18, 20, -18, 1, 19, -7, -15, -21, 38, 70, 49, 24, -29, 15, 37, 21, 16, 18, 6, 9, 10, -24, -32, -50, -8, -60, 13, 48, -2, 13, -18, -19, -8, 19, 4, -20, 57, 22, 36, 19, 34, 33, 65, 41, 26, 8, -16, -19, -21, -39, -56, -37, -52, -88, -30, 10, 20, -2, 7, 0, -20, -5, -7, -21, 13, -7, 16, 17, 48, 39, 22, 45, 7, -40, -48, -36, -54, -83, -82, -56, -63, -79, -46, -23, 8, -30, 4, 16, 6, 4, 17, -82, -17, 14, 9, 43, 54, 41, 38, 34, 19, -55, -77, -56, -105, -70, -90, -69, -103, -64, -66, -15, 8, 11, 2, -10, 15, 21, -33, -81, -16, -10, 29, 59, 33, 61, 71, 37, 31, -18, -7, -24, -32, -34, -38, -15, -99, -29, -27, -7, -5, -4, -14, -17, 2, -19, 4, -43, 4, -11, 23, 11, 10, 47, 45, 45, 41, 25, 73, 8, 27, 27, -14, -19, -17, 2, 14, -21, 16, -13, 9, -15, 17, 14, -15, -37, -30, -27, -22, -39, -22, 1, -4, 8, 11, 42, -4, 29, 53, 34, -4, -8, -16, 13, 56, 36, 17, 8, 7, -12, -2, -18, -41, -28, -2, -40, -22, -16, -18, 22, -10, 7, 10, 19, -4, 10, 22, 19, -3, 12, 19, 23, 55, 23, 48, -9, 15, 14, 13, -19, -18, 22, 14, -10, -12, 5, 4, 19, -33, -33, 0, -14, -11, -7, -8, 6, 1, 27, -22, 28, 58, 50, 49, 27, -17, 1, -16, -12, 52, 49, 31, 16, -5, -4, -13, 26, 2, -3, 19, -17, -13, 15, 0, 24, 61, 29, -11, 1, 51, 38, 37, -9, 19, 8, -14, -5, 47, 43, 34, 31, 10, 33, 48, 36, 24, 48, 24, 34, 26, 34, 5, 67, 44, 45, 49, 13, 33, 31, 43, -16, -19, -19, 7, 0, 41, 34, 43, 1, 11, 37, 29, 31, 4, 48, 47, 32, 86, 67, 60, 31, 32, 28, 49, 24, 21, 19, 55, -23, -19, 17, -5, 7, 80, 49, 31, 2, -15, 16, 18, 30, 31, 14, 27, 35, 42, 50, 59, 57, 52, 41, 45, 16, 9, 37, 33, -1, -15, 2, -10, 10, 29, 42, 26, -7, 20, 14, 48, 27, 35, 16, 23, 41, 25, 29, 26, 78, 69, 38, 54, 39, 35, 39, 22, 6, -7, -4, -8, 10, 23, 7, 22, 27, 39, 22, 26, 48, 25, 27, 38, 28, 14, 24, 12, 55, 81, 27, 65, 49, 62, 28, 37, 16, 7, 6, -3, -18, -7, 18, 44, 2, 32, -1, 54, 42, 28, 13, -12, 23, 10, 10, -17, 20, 38, 47, 30, 12, 24, 41, 17, 24, -15, 18, -2, 18, -6, -25, -33, 21, 20, -7, 20, 24, 7, 2, 9, -15, 11, 13, 16, 33, 7, 49, 6, 12, -1, -7, 16, -2, 18, -19, -16, -13, 39, -12, 14, 20, 14, 0, 22, 1, 12, -11, 23, 24, 14, 18, 0, 13, 25, 32, -1, 11, 20, 29, -10, 39, -14, -18, 16, 5, 41, 63, -14, 2, -11, -9, -17, 1, -14, -27, -39, -32, 2, 9, 16, -10, 9, 12, 29, 21, 30, 13, 0, 40, 2, 3, 20, 15, 1, 41, 47, 71, 55, 68, 57, 47, 4, 10, 10, -13, 9, 41, 52, 50, 65, 22, 47, 14, 26, 53, 33, 0),
  72 => (9, 13, 6, 4, 17, 0, -5, -1, -10, -3, -14, 0, -9, -16, 10, -2, -33, -31, -18, -31, 2, -10, 17, -17, 15, 14, 20, -15, -14, -11, -17, -20, -3, -2, -20, -18, -7, -1, -7, -19, -25, -36, -15, -12, 3, -22, -22, -12, -10, -21, -19, 12, 13, -9, -1, -6, -8, 8, 19, -1, 5, 3, 4, 13, 13, -21, -27, -14, -34, -16, -10, 9, -4, -24, -11, -56, -25, -14, -34, -65, -6, -1, 16, -14, -16, 8, 5, -17, 18, 1, 19, 16, -5, -19, -32, -48, -19, 19, 30, -2, -48, -37, -39, -21, -19, 5, 7, -51, -38, -41, -17, 19, -11, 12, 7, 4, 19, 19, -10, 5, -15, -36, -78, -21, -8, 56, 8, 3, 7, -11, -15, -8, -24, -43, -41, 17, -7, -32, 1, -9, -19, -20, -3, -12, -14, 12, 4, -15, -37, -27, -60, -22, -10, -26, -6, -32, -15, -19, -15, -15, -29, -24, -18, 33, 24, -13, 0, 4, 9, 16, 19, -10, -8, -8, 4, -78, -8, -36, -7, -9, -26, -19, -30, -62, 5, -4, -42, -14, 0, 2, 5, 43, 41, 10, -12, 4, 10, 15, -14, -5, -12, 20, -30, -39, -46, -18, -6, 15, 1, 13, -40, -33, -33, -22, -4, 9, -6, 3, 3, 35, 7, 9, 5, 19, 12, -17, 5, -10, 10, 8, -42, -12, -19, -11, -8, 0, -34, -36, -49, -40, -47, -31, -20, 14, 6, 19, 59, 45, 55, 18, -16, -10, 17, -13, -17, -5, -8, 18, -56, -4, 0, -5, -27, -18, -28, -32, -29, -8, -22, -20, 20, 42, -7, 56, 60, 66, -2, -22, 7, 12, -2, -7, -5, 18, -8, 16, -17, 48, 32, 42, 21, 37, 29, 11, 0, -27, 2, 7, 7, 50, 20, 62, 40, 14, 25, -8, 10, -26, 15, 7, 9, -11, 9, 31, 91, 65, 26, 51, 19, 21, -7, -6, -20, 0, 16, 21, 6, 44, 45, 51, 49, 7, 15, -4, -6, -39, -6, 20, 1, -15, 12, 22, 77, 51, 1, 63, 20, 15, -18, 11, 20, 16, -2, 21, 19, 33, 76, 0, 8, 13, 17, -13, -1, -63, 19, -17, -15, 19, -38, 10, 76, 15, 36, 56, 20, 17, 22, 28, 46, 20, 24, 21, 26, 53, 64, -17, 0, 5, 37, 21, -11, -31, 19, 10, -19, 13, -64, 16, 54, 35, 47, 23, -26, 17, 23, 34, 26, 55, 57, 39, 14, 11, 29, -2, 2, -9, 2, -4, -28, -23, 1, 6, 8, -9, -26, 0, 44, 42, 15, -20, 16, 34, 15, 2, -1, 34, 40, 34, 22, 1, -9, 8, 16, 22, -11, -19, -50, -2, -8, 12, -1, -7, -19, 37, 22, 39, 21, 2, 11, -11, -13, -2, -1, -5, -33, -12, -29, -23, -38, -16, -2, -20, -19, -51, 16, 10, 15, -12, -1, 16, -19, 16, -22, -3, 4, -24, -46, -12, 8, -22, -7, -57, -20, -54, -84, -54, -54, -58, -65, -79, -36, -37, 2, 59, 12, -8, -12, -16, -27, -48, -25, -1, -16, -17, -34, -61, -53, -35, -53, -84, -70, -56, -59, -40, -38, -81, -93, -77, -74, -57, -49, 35, 16, 7, 5, -11, -56, -49, -13, -7, -5, 16, -1, -38, -53, -49, -74, -67, -51, -84, -47, -12, -44, -46, -60, -60, -62, -66, -49, 17, -3, -3, -16, 19, -53, -65, -14, 6, -9, -25, -25, -83, -34, -22, -44, -54, -53, -72, -20, -49, 4, -18, -66, -36, -82, -52, -22, 1, 10, -4, -13, -6, -17, -47, -32, -5, -14, -71, -40, -41, -17, -2, -40, -57, -30, -9, -35, -60, -12, -30, -36, -24, -48, -55, -55, 4, 10, 18, 12, -18, -59, -37, 2, 7, 3, 6, -36, -19, -31, -54, -33, -48, -74, -46, -48, -68, -20, 9, -38, -66, -32, -44, -29, -17, -16, -13, 16, -1, -23, -53, -18, 39, 33, 7, 0, -8, -51, -55, -65, -37, -49, -67, -30, -43, -63, -10, -12, -33, -25, -33, -1, -22, -19, -2, 14, 0, -37, -56, -21, -8, 2, -14, -45, -48, -44, -61, -26, -32, -14, -58, -47, -26, -58, -29, -4, -30, -3, -13, 3, -1, 4, 17, -20, -7, -18, -22, 16, 21, 29, 16, -25, -44, -4, -25, -21, -29, -2, -38, -17, -18, 13, -16, 6, 9, -13, 15, -19, -31, -1, -19, -11, -13, -15, -26, 2, 3, 2, 26, -29, -41, -53, -34, -1, -47, -20, -26, -12, 8, -25, -29, 11, 1, -4, 4, -5, -19, -10, 12, -6, 17, -8, -2, 17, 20, 14, 5, 13, 2, -4, -6, -22, -20, 3, -8, 0, -12, 0, 8, -15, -15, -6, 5, 6, -14),
  73 => (-1, 13, 6, 4, -15, -20, -16, -6, 1, -4, -6, 9, 18, 12, 19, 25, 81, 60, 69, 35, 45, -2, 15, -1, 4, 9, -5, -13, -5, -13, 15, 6, -14, -14, 2, -3, -11, 14, 9, -19, -24, -24, -32, -2, 24, 40, -5, 2, 22, 20, 14, -11, -17, -12, 14, -8, 17, -16, -11, -4, -1, 15, 18, 7, 8, -7, -3, -39, -74, -66, -32, 10, 56, 38, 36, -3, -17, -10, 24, 21, -18, -24, -8, -6, 3, -11, -13, -16, 8, -12, 11, -5, -22, -51, -31, -21, 7, 1, 43, 70, 41, 30, -14, -7, -24, -47, -31, 6, 5, 14, 20, -4, 15, 11, -6, -6, 10, 9, 21, -3, -25, 4, -41, -27, 10, -9, 1, 46, 41, 37, 30, 14, 31, 17, 8, 24, 42, 1, 1, 17, -4, -20, 19, 19, -8, -1, -28, -13, -9, 0, 10, -6, 7, 28, 41, 53, 61, 56, 65, 62, 34, 58, 39, 12, -14, -5, 19, -3, -3, 16, -7, 15, -14, 16, -20, -4, -41, 26, 42, 18, 18, 51, 67, 76, 87, 63, 73, 80, 46, 97, 43, 26, 44, -36, -29, -7, -18, 12, 13, -20, -19, -19, 26, 34, -4, 26, 16, 22, 39, 59, 84, 113, 106, 83, 87, 58, 45, 67, 64, 45, 37, -66, 13, 1, 6, -4, -15, -12, 4, 20, 30, 53, 39, 47, 60, 43, 47, 62, 84, 84, 54, 48, 16, 46, 45, 64, 64, 50, -4, -7, -5, 31, 13, -18, -14, -17, -18, -17, 30, 32, 49, 92, 51, 8, -16, -17, -33, -52, -49, -43, 13, 2, 14, 8, 8, -1, -28, 13, -16, 34, 1, -16, 11, 20, 4, -8, 59, 44, 49, 36, -7, -60, -58, -37, -33, -18, -8, -56, -15, -2, -8, 6, -18, 0, -14, -5, -11, 20, -6, 9, -4, -5, -11, -45, 16, -14, 25, 12, -13, -5, -23, -21, -22, -9, -13, -69, -47, -30, -28, -5, 4, -18, -39, -44, -35, 28, -10, 17, 1, 8, -8, -78, 9, 5, 25, 23, -11, -17, -10, -23, -25, 13, 19, 1, -2, -18, -14, -10, -27, -56, -69, -46, -74, -18, -9, 10, -11, -13, -19, 1, -26, -25, -24, -6, 11, 19, -7, -9, -5, 30, 64, 10, 14, -11, -10, -21, -38, -54, -36, -48, -54, -5, -21, -18, 19, -15, 11, 33, -33, -64, -38, -18, 8, 6, 11, -17, -22, -17, -3, -8, -20, -9, -28, -4, 24, -17, -36, -33, -78, -14, -7, -19, 18, -3, 11, 25, 12, -68, -38, -24, -61, -31, -4, 17, -20, -19, -25, -21, -66, -23, -16, 8, -9, -6, 7, -31, -72, -6, 9, -11, 2, 4, -52, -13, -6, -46, 9, -16, -23, -16, -3, 12, -7, -9, -39, -32, -5, -24, -23, -7, 10, 3, -27, -27, -35, 2, 5, 6, -14, -2, -54, 24, -30, -20, 27, -3, -15, -2, -17, -1, -34, -32, -65, -50, -10, -29, 9, -1, -5, 5, -34, -42, -31, 21, -2, 9, -18, -11, 2, 13, -25, 0, 9, 25, 25, 20, 12, -14, -46, -5, -31, -27, 18, 0, 7, -5, -11, 48, 15, -28, -30, 0, -18, 1, 8, -6, -15, 7, 16, 7, 9, 13, 14, -14, 15, 0, -9, -7, -43, 4, 21, -12, 15, 5, 7, 15, 26, -23, -35, 29, 19, 8, -15, 6, -33, 15, -17, 5, 17, -4, -10, 0, -4, -7, 6, 11, -42, -30, 6, -23, 6, 21, 19, 17, 29, 26, 1, 19, -1, -12, -13, 3, -13, 16, 31, -6, 4, -31, 1, -8, -15, -47, -33, -22, -47, -40, -6, -4, -2, -11, -14, -27, 36, -11, -33, 9, 10, -7, -7, -11, -58, 34, 70, 8, -15, -31, 14, 10, -6, -9, -9, -7, -47, -10, -15, -5, 4, -11, -32, 3, 19, 41, -22, 24, 3, 0, -4, -13, -46, -18, 61, 53, 22, -6, 10, 17, 14, -17, 28, -9, -32, -13, -25, -25, -35, -50, -10, -4, 35, 1, -4, -17, 0, 4, -2, 2, -31, 10, 2, 3, 43, 3, 26, 23, 21, 2, 20, -2, -23, -27, -27, -36, 5, 8, 0, 1, 14, 19, 32, 2, -7, 11, 0, -14, -8, -27, -13, -5, -20, 2, 23, 27, -6, -3, 18, -1, -19, 27, -2, 23, -13, -3, -28, 27, -1, 21, 13, -6, 2, 18, 5, 14, -12, -12, -43, -24, -25, 0, 1, -17, -20, -10, 5, 17, -18, 24, 24, 18, 24, 8, -27, 36, 18, 13, -9, -13, 3, -16, -3, -3, -4, -8, -9, -33, -33, -31, -46, -30, 11, 30, 23, 8, -30, -35, 8, 4, -2, -4, -8, 14, -14, 5, -3, -5),
  74 => (-9, -4, 14, -18, -10, -1, -9, 2, -17, -18, -1, 18, 18, -6, -1, -2, 8, 18, 29, 48, 26, -5, 7, -19, -11, -6, -9, -18, 6, -8, -13, -19, 14, -14, -1, 9, -8, 20, -1, -20, -10, 8, 14, -17, 11, 12, 22, 44, 26, 16, 13, 20, 16, 3, -12, 17, -18, 11, -8, -19, 20, 3, 14, 20, 11, 0, -14, -2, -11, 8, 12, 45, 35, 13, -3, -32, 10, -9, 32, -19, -27, -17, -16, 17, -7, 8, -17, 11, 10, 4, 16, 14, -23, 0, 14, 3, -12, -3, -26, -59, -21, -12, -26, -7, -18, -10, 10, -22, -2, 6, -21, -18, -12, -13, 17, -6, -6, 11, -14, 9, 14, 32, 4, -23, -31, -45, -90, -45, -33, 31, 43, 12, 29, 18, 2, -37, 3, -6, -3, 9, 6, 1, 5, -16, -16, -17, 2, -6, 42, 18, 5, -59, -68, -96, -56, -40, 2, 68, 15, 30, -2, -24, -38, -42, -27, -22, -14, -2, -18, 20, 2, 5, 4, -13, 14, 13, -1, -26, -5, -37, -79, -110, -66, -11, 14, 66, 22, 5, -15, -31, -43, -70, -25, -13, -11, -17, -10, -10, -17, -11, 17, 18, 47, 27, -3, -19, -21, -30, -113, -112, -52, -16, 26, 51, 6, 17, -22, -19, -66, -50, -48, -41, -10, -20, -15, 19, 1, -18, 8, -16, 43, 4, 2, 7, -18, -34, -110, -87, -70, -6, 15, 43, 8, -20, -32, -35, -58, -54, -70, -27, 3, -19, 18, 2, -4, 14, -14, 14, 6, 0, 18, 11, 8, -15, -36, -69, -44, 8, 14, 53, 6, -33, -14, -42, -36, -39, -18, -37, -34, 9, -20, 16, -6, -1, 3, 12, -32, 58, 10, -24, 11, -37, -39, -79, -66, -14, 6, 21, -17, -27, -37, -44, -33, -16, -17, -50, -17, -1, -8, -5, -15, 16, 7, -24, 26, 78, 25, -34, -28, -42, -82, -62, -42, -37, 2, 15, -26, -27, -27, -55, -1, 22, -7, -15, -32, -32, 6, -17, 0, 6, -9, -5, 50, 36, -13, -7, -2, -36, -46, -48, -19, -9, 13, 20, 2, -2, 15, 4, -22, 10, -10, -38, -21, -11, -11, -8, 20, 8, 17, 32, 61, 6, -5, -15, -27, -20, -40, -56, -6, 9, 30, 17, 30, 17, -10, 3, -7, 0, 27, 5, -24, -48, 7, 11, 7, -4, 1, 11, 61, 7, -5, -13, -69, -19, -51, 1, -21, 13, 9, 14, 35, -16, -28, -8, -13, -19, -4, 8, -6, -19, 7, 11, -14, -16, -1, 26, 1, 19, -8, -5, -18, -27, -26, -2, 14, 14, -11, 20, 15, 46, 36, 19, -26, -5, -21, -10, -11, -8, -8, -3, 12, 16, 30, 45, 6, 7, 16, -18, -38, -9, -38, -12, 36, 17, -12, 10, 11, -17, -14, 12, -39, -2, -4, -31, -2, -45, 6, 21, -6, -1, 39, 33, 8, 13, -23, -41, -78, -29, -63, -26, 3, 1, 10, -27, -26, -4, 4, 1, -17, 10, -12, -16, -1, -16, -20, -4, 17, -10, 74, 55, 20, -2, -9, -23, -57, -109, -73, -25, 9, -21, 24, -4, -30, 5, 26, 5, 12, -1, 0, -2, -2, -36, 3, 1, 14, -7, 21, 9, 34, 5, -46, -4, -21, -46, -63, -11, -4, -1, 1, 20, -16, 2, 5, 14, -14, 11, 9, -36, -36, -58, -16, 9, -19, 12, 10, -7, 31, 18, -2, 28, -7, -2, -66, 8, -4, -3, 23, 32, 22, 1, 28, 6, -23, -29, 6, -38, -6, -12, 12, 16, -20, -19, -5, 11, 24, -24, -8, 21, 40, -14, 1, 29, 40, 28, 37, 16, 23, 43, 28, 20, 23, -17, -2, -25, -13, -18, -8, 9, -17, -3, -19, 10, 6, -3, 11, -9, 8, -2, -2, 72, 58, 75, 60, 48, 3, -36, 21, 4, 10, -18, -18, -8, 10, 21, -11, -13, 3, 13, 17, -7, -20, -18, 11, 53, 2, 0, 37, 37, 29, 49, -4, -4, 8, -18, -11, -17, -22, -15, 3, 8, 8, 26, 21, -6, 17, -17, -1, 11, -12, -22, -31, 8, 13, -3, 38, 34, 63, 41, -4, 4, 39, -9, -10, 7, 9, 1, -33, 1, 18, 41, -7, -3, 8, -8, -19, 26, 20, -32, -35, -32, -25, -14, -6, -7, -22, 46, -11, -17, 13, -19, -3, -1, -30, 0, -28, -16, 3, -21, -18, 1, 11, 19, 17, -18, 13, -10, 17, -11, -34, -43, -54, -29, -41, 8, -14, -7, -5, -26, -6, 4, -38, 7, 35, 9, -13, -26, -9, 19, 18, -2, -1, 18, -6, 3, -4, -18, -32, -9, -16, -22, -5, -31, -21, -5, 30, 23, 14, -22, -37, -45, -25, -9, -48, -41),
  75 => (8, -8, -4, -18, 19, -13, -5, -2, -8, -7, 15, -5, 17, -9, -21, -32, -24, -10, 1, -22, 7, 7, -12, -11, 13, -10, -7, 20, 4, 19, 15, -16, -14, -1, 19, 11, -3, -6, -4, 5, -38, -9, -34, -42, -74, -31, 5, -19, -2, -20, -4, 3, 2, 9, 20, -6, 14, 0, 9, -8, 18, -11, 10, -13, -8, -16, 1, -26, -33, -69, -72, -13, 7, 43, 40, -14, -29, -19, -39, -30, -19, 15, 18, 6, 15, 3, -18, 11, -16, 8, -15, -16, -20, 44, 39, 17, -33, -64, -2, 50, 26, 36, 15, -8, -38, -50, -39, -14, -16, 7, 10, 8, -1, -2, -16, 11, -8, -11, -6, -23, 61, 39, 28, -12, -25, -9, 45, 12, 13, 15, 9, -20, -5, -72, -36, -13, 2, 11, 9, 5, 8, 7, -17, 8, -8, -6, 11, 2, -56, -40, -61, -36, -7, -23, 21, 53, 20, 7, -3, -7, -8, -48, -27, -15, -35, -20, 0, -3, -4, -11, 4, -16, 7, 15, -17, -2, -56, -44, -66, -63, -15, -26, 16, 3, 32, 6, 1, -8, 6, -18, 20, -2, -32, -18, -20, -5, 10, -10, -12, -3, -4, -6, 22, -18, -59, -65, -86, -38, -41, 0, -4, -3, 3, 7, 20, -2, -16, -8, -11, 32, -15, 7, -14, 9, -11, -7, -9, 7, -7, 9, 0, -25, -63, -108, -66, -82, -45, -30, -13, 7, -16, -11, -37, -23, -4, 3, 45, 14, 9, -15, 39, 2, -1, -4, -2, 12, 0, 11, -28, -34, -77, -100, -50, -14, -28, -33, -42, -27, -14, -14, -5, -23, 6, 38, 19, -1, 4, 31, 33, 18, -18, -14, -4, -8, 3, -28, -30, -63, -58, -38, -17, 16, -6, -15, 9, 7, -32, -34, -25, -5, 0, -7, 24, 23, 6, 0, -22, 1, 11, 0, 20, -2, -16, 17, -33, -48, -39, -21, 24, 45, 38, 44, 31, -14, -57, -49, -14, -23, -10, -3, 13, 31, 23, 19, -7, 8, 3, 15, -4, 13, -8, -5, -10, 0, 6, -4, 59, 60, 70, 58, -8, -8, -35, -27, -39, -2, 5, -10, 19, 16, 9, 4, -51, 29, -7, 2, -12, 14, 12, 16, 29, 32, 10, 14, 68, 89, 57, 67, 30, -7, -17, -12, -11, 5, 5, 27, 22, 16, 5, -38, -52, -35, -7, -5, 4, 12, 6, -14, 18, 7, -22, 13, 46, 66, 47, 60, 50, -6, -25, -25, 6, 6, -1, 21, 13, 19, 6, -43, -8, -8, -3, -11, -4, 3, -44, -40, -34, -45, -53, -6, 49, 32, 40, 50, 80, 30, -3, -2, -8, 9, 1, 26, 16, 5, -10, -37, -48, 28, 6, -13, -18, -15, 40, -38, -30, -50, -46, -34, 12, 29, 23, 36, 66, 37, 5, -3, -15, 12, 14, -2, 0, -11, -12, -43, -33, 22, -8, -16, 17, 8, -16, -20, -28, -49, -75, -47, 18, 14, 36, 1, 37, 12, 2, 14, -5, 10, 44, 10, -3, -18, -10, -5, -12, 5, -2, -7, 9, 17, -24, 6, -47, -67, -100, -60, -46, 13, 15, 3, -13, -5, 0, 26, 24, 20, 39, 3, 27, 16, -21, -19, 6, 18, -11, 8, 12, 8, -7, -18, -31, -57, -93, -56, -55, -27, 9, 24, -8, -10, -37, -1, -10, -29, 14, 31, 32, 53, 58, 12, 2, 30, -4, -2, 6, 17, -17, -18, -75, -69, -106, -41, -89, -65, -30, 37, -33, -16, 1, 14, 19, -4, 26, 8, -35, 23, 16, -13, -3, 41, 4, -16, 2, 2, -8, -32, -26, -20, -39, -43, -57, -133, -58, 6, -29, -20, 1, -27, -12, -3, -9, -16, -64, -5, 17, 12, 3, -2, 10, 13, 9, 16, -19, -24, -19, -35, -13, -7, -48, -124, -114, -64, -28, -10, -13, -4, 26, 7, -2, -41, -44, -56, 13, 28, -11, 14, 20, 0, 1, -9, 0, -23, -8, -7, 10, -18, -50, -114, -49, -56, -78, -48, -33, -23, -40, -10, -68, -72, -68, -45, -6, 15, -30, 27, 7, 20, 2, 4, -2, 5, 10, 14, 27, 20, -34, -99, -87, -60, -49, -70, -80, -58, -75, -33, -89, -79, -49, -51, -61, -13, -31, -11, -14, -14, 2, -12, -3, 16, 20, -15, 2, 31, -2, -53, -37, -32, -53, -37, -35, -39, -62, -55, -34, -53, -14, -75, -59, -68, -13, 0, 5, 10, -10, 13, 22, 0, 11, 15, -6, -36, -24, -15, -18, -32, -48, -38, -52, -59, -31, -50, -22, -23, 5, -55, -23, -56, -25, 5, 4, -21, 11, 20, -11, 19, -19, 12, -4, -1, -11, -20, -13, -10, -40, -24, -15, -15, -26, -29, -48, -41, 10, -30, -63, -32, -5, 1),
  76 => (-6, 0, -10, -16, 15, -4, -14, -3, -17, -2, 2, -13, 10, -15, 26, -21, -20, -28, -47, -84, -28, -9, -43, -1, 19, -2, -13, -7, 7, 10, -19, 2, -6, -2, 8, 3, 6, -12, 29, -11, 16, 47, 65, 56, 44, 19, 1, 19, -26, 14, 34, -17, -18, 19, 17, -18, -4, -10, 3, -15, -5, -5, 11, -18, 11, 27, 26, 76, 79, 75, 80, 41, 47, 47, 61, 39, 33, 17, 19, -16, -77, -27, -17, 1, -2, 14, 11, -1, 6, 2, 0, 2, 56, 62, 46, 36, 57, 71, 46, 1, 0, 13, 23, 34, 27, 27, 6, 31, 2, -23, -4, -14, 15, 14, -11, -3, -20, 13, 0, 21, 58, -20, 30, 29, 7, 26, 30, 15, 15, -9, 38, 7, 0, 6, -5, 0, -20, -26, 7, 7, -18, -4, -11, 9, 6, 5, 36, 52, 19, 5, 25, 37, 46, 52, 33, 50, 29, 17, -6, 5, 11, 11, 25, 3, -5, 9, -12, -15, -3, 9, -19, -10, -20, -7, 13, 17, 10, 26, 60, 22, 51, 35, 50, 32, 16, 4, 14, 17, 26, 20, -7, -8, 30, 4, 15, -17, -16, -7, 1, 16, -4, -17, 37, 44, 34, 68, 35, 31, 14, 32, 24, 31, 33, 13, 19, 32, 25, 32, 24, 17, 6, -15, 25, 4, 6, -4, 7, -12, -16, -16, 14, 56, 51, 71, 30, 7, -12, 15, 16, 53, 18, 22, 31, 19, 30, 4, -1, -10, -8, 13, -20, 2, -20, -8, -1, 5, -17, 0, 11, 66, 40, 65, 15, -9, 12, 13, 54, 31, 5, 31, 36, 23, 37, 25, 38, 16, 4, -3, -7, -34, -13, -11, -7, -9, 16, -15, 22, 51, 39, 24, 6, 46, 49, 40, 55, 47, 8, 68, 48, 44, 75, 42, 5, 16, 7, 5, 20, -52, -5, 3, 14, 11, 0, -52, 16, 14, 14, -4, -7, -2, 30, 17, 15, 39, 34, 29, -5, 29, 16, 32, 8, 3, 28, 24, 24, 12, -13, -7, 21, 3, 24, -69, 53, 9, 27, 28, 11, -8, 4, -17, 8, 5, 20, -5, 2, 12, -19, -13, -3, 25, 72, 63, 43, 18, 12, 9, -7, 6, -37, -76, 5, 19, 36, 45, 23, -15, -13, -24, -2, 28, 35, -4, 18, 19, -31, -28, 35, 14, 47, 51, 30, 55, -2, -9, 8, -16, -43, -36, -9, 14, 64, 50, 61, 43, 19, 49, 80, 41, 51, 12, 22, 51, -8, -13, -14, -1, 35, 23, 22, -3, -5, 20, -10, 10, -62, -32, 11, 12, 54, 56, 59, 65, 61, 64, 77, 102, 68, 62, 40, 54, 25, 21, 23, 15, 39, 21, -12, 11, -15, -8, 4, -3, -20, -30, 42, 99, 105, 60, 66, 61, 94, 64, 103, 74, 47, 29, 50, 52, 30, 36, 43, 13, 22, 9, -51, 8, 19, 12, -10, 8, -14, 35, 65, 103, 72, 32, 48, 19, 60, 48, 42, 19, 38, 35, 40, 8, 22, 28, 39, 30, 21, 17, 14, 14, -7, -10, -14, -16, 8, 32, 53, 40, 29, 13, 6, 1, -7, -25, -12, 39, 1, 25, 46, 14, -2, 16, 5, 20, 29, 12, 27, -30, -14, 10, 15, 14, -3, 30, 27, 1, 38, 35, -16, 0, -39, -29, -12, 18, -17, 11, 30, -4, 5, 28, 25, 30, 27, 16, 36, -24, 12, 17, 0, 12, -23, 26, 8, 11, -2, -18, 9, -7, -9, -16, -4, 0, -23, -37, -22, -41, 7, 43, 43, 21, 35, 41, 38, -29, 12, 8, -5, -4, -58, 1, 42, 6, 25, -3, 42, 7, 22, 12, 42, 39, 17, -14, 13, 20, 39, 64, 40, 46, 56, 21, 37, -44, 20, 8, 15, 14, -63, -11, 16, 9, 9, 2, 28, 11, 21, 23, 30, 29, 7, 26, 27, 4, 28, 49, 36, 35, 34, 36, 19, -28, 16, 1, 5, 11, -56, -18, 18, 25, 27, 42, 2, -33, -2, 17, 7, 4, 28, 33, 6, 23, 56, 67, 58, 28, 37, 20, 30, -17, -14, 16, -10, 1, -40, -36, 9, 34, 13, 41, 32, 34, 31, 6, -4, 1, 22, 37, 8, 24, 28, 67, 21, 29, 54, 33, 52, -43, 14, -7, -10, -13, -66, -37, 18, 26, 0, 3, 41, 33, 25, 31, -4, -13, 14, 19, 30, 12, 42, 31, -2, 7, 42, 23, -15, -50, -3, 20, 7, -4, -7, -6, 23, 4, 7, 9, 31, 29, 12, 18, 16, -20, -6, 29, 33, 46, 19, 14, 20, -24, 12, -1, -48, -44, 5, -12, -11, -12, 9, 54, 75, 73, 31, 23, 46, 53, 22, -5, 34, -3, 23, 71, 40, -30, 18, -15, -16, -20, -9, -18, -75, -46),
  77 => (-18, 17, 4, -12, -18, -15, 14, 0, -8, 13, 2, -5, 3, 6, 5, 25, 38, 56, 42, 29, 27, -22, -3, 6, 1, -10, -19, -14, -19, 4, 3, -7, -15, -17, -20, 12, 10, 9, 5, 21, 32, -4, -34, 5, 33, 21, 17, 16, -7, -14, -28, -9, 13, -14, -7, 19, -19, -3, 16, -8, -7, 19, 7, 10, 6, -25, -29, -18, -44, -13, 6, -13, -17, -16, -10, 4, -1, -10, -13, 7, 36, -1, -18, 1, 2, 0, -3, -8, 18, 4, -5, 5, 2, 23, -19, -15, 30, 5, 24, -7, 33, -21, -1, -27, 17, -14, 15, 31, 53, 21, 5, -20, 0, -11, 8, 11, -9, 13, 5, -10, -15, -8, -25, 12, 11, 6, 17, 25, 42, 23, 1, -21, 17, -7, 7, -37, 10, 13, 7, -10, -2, 16, -9, -2, -7, -10, -34, -3, -59, -13, -1, -15, 3, 31, -15, -23, 1, -17, -21, -3, 26, 5, 3, -13, 0, -3, -11, -18, -11, 17, -15, 5, 15, -15, -30, -42, -39, 2, -7, -6, 8, 14, 0, -11, 8, 5, 4, -22, 15, 9, -4, 18, 3, 16, 6, -7, -14, 10, -9, 11, 8, -10, -13, -2, -10, -35, 21, 10, -17, 10, -14, 3, 1, 6, 9, 9, -4, 20, 6, 25, -6, 11, -1, -9, -3, -2, -16, -16, -9, 7, -45, 30, -18, -63, -4, -1, -3, 10, 2, -31, -32, -7, 14, 7, -6, -1, -9, -4, -5, -4, 23, -15, -6, 0, 20, -5, -9, -16, 41, 25, -15, -31, 7, -17, 32, 26, 3, -55, 10, 36, 32, 24, -9, 23, 17, -42, -1, 11, -1, 5, 6, -8, 11, -18, -3, 27, 63, 28, -1, 12, 3, 3, 38, -1, -43, -71, -25, 26, 10, 20, -12, -15, -4, -38, -28, -7, -26, 16, 10, -9, -20, 16, -18, 0, 68, 39, 9, 20, -3, -19, 44, -5, -71, -69, -10, 34, 2, 7, 5, -19, -19, -26, -20, 4, -26, -15, -2, -9, -18, -9, -3, -36, 24, 16, -6, 19, 15, 13, 42, -15, -68, -81, -6, 34, 13, 8, 33, -4, -55, -43, -24, -31, 7, -4, 12, 20, -8, -5, -22, -11, 38, -55, -47, 13, 12, 17, 68, -24, -70, -96, -27, 40, 4, 25, 15, -20, -36, -20, -49, -33, 21, 10, 0, 3, 15, 9, -6, 73, 21, -43, -38, 46, 19, 17, 19, -43, -76, -112, -13, 44, 17, 21, 28, -20, -38, -38, -45, -9, 2, -20, -20, -4, 4, 13, 47, 50, -24, -61, -56, 27, -5, 13, 21, -30, -77, -93, -10, 29, 13, 26, 6, -20, -32, -35, -31, -35, -1, -37, 18, -1, -6, 10, 5, 14, -68, -68, -17, 39, 15, 17, 48, -44, -114, -118, 22, 22, 0, 54, 29, -22, -41, -49, -56, -45, -29, -40, -6, -16, -3, -16, 13, -36, -84, -84, -10, 25, 37, 30, 51, -6, -113, -85, 26, 46, 11, 30, 19, -47, -60, -67, -50, -31, -7, -36, -9, 0, 13, 14, -5, -60, -91, -42, -30, 6, 18, -7, 10, -17, -94, -96, 24, 27, 12, 43, 12, -14, -47, -42, -46, -34, -27, -17, 10, -17, 2, 17, -11, 5, -49, -66, 20, 34, 38, -17, 10, -37, -102, -65, 20, 40, 20, 20, 6, -23, -24, -69, -67, -32, -10, -19, -9, -17, 2, 9, 18, -10, -48, -3, -12, 24, -3, 14, -10, -5, -76, -46, -5, 40, 32, 30, 2, -27, -34, -59, -32, -6, -17, 18, 8, -13, 15, 4, -7, -19, -31, -24, 27, 6, -1, -10, -9, -44, -81, -50, 7, -4, 24, 55, 1, -27, -13, -48, -35, -16, 16, 7, -18, 16, -12, -18, -28, -13, 22, 51, 14, 10, -21, -5, -16, -23, -75, -29, 24, 36, 33, 52, 7, -23, 9, 7, -45, 4, -5, 33, -14, 19, -17, -11, 14, -5, 7, 38, 20, -12, -11, -21, -11, -52, -46, -35, 33, 29, 39, 25, 30, -48, -47, -33, -38, -17, -6, -18, 16, 16, -9, 9, 0, 23, 11, 3, 16, 8, -17, -59, -53, -44, -35, 17, 25, 23, 36, 47, -20, -21, -22, -29, -11, -28, -30, 18, -16, -15, 2, 7, -12, 14, 7, -8, 24, -3, -44, -62, -64, -76, -33, 49, 26, 12, 36, 17, -20, -44, -13, -43, -21, -4, -19, -1, 9, 18, -7, 20, 18, 6, -26, -12, -2, -6, -43, 3, -61, -52, -13, 16, 27, 23, -2, 14, -28, -2, -18, -46, -35, -23, -3, 11, 5, -18, -19, -4, -17, -8, 4, 14, -25, -12, -19, -23, 23, -35, -14, -1, 37, 17, 39, -12, 3, 33, -17, -45, -45, -17, -39, 7),
  78 => (2, -18, -13, -18, -10, 9, 20, 11, 4, -1, -14, -7, 3, 17, -10, -58, -56, -6, 15, -16, -65, -43, -5, -19, -5, 13, -18, 15, -4, -14, 20, 20, 19, 18, -19, -15, 7, 10, -4, 52, 74, 20, 39, -17, 2, -14, -7, 26, -2, -11, 33, -31, -40, -15, -1, 19, -5, 16, 5, 6, -20, -3, 14, 4, -6, 23, 62, 54, -13, -14, 27, 10, -17, 15, 13, 3, -8, 12, -8, -11, -22, -22, -17, -19, 12, 19, 12, 18, 16, -5, 21, 11, 49, 87, 72, 45, 57, 81, 26, 15, 9, -8, 25, 6, -14, -16, -21, -15, -18, 26, 14, -8, 2, -20, -5, 15, 15, 7, -10, 46, 54, 52, 73, 72, 15, 60, 40, 40, 84, 29, 35, -12, -31, -5, -17, -12, -32, -21, 4, -2, -10, 10, 5, -4, -19, -19, 35, 80, 52, 5, -3, 27, 65, 49, 47, 54, 58, 24, -21, -16, -29, 13, 13, 9, 14, -18, 2, 9, 15, 16, 17, -15, 18, 6, 59, 124, 20, 31, 22, 47, 54, 58, 59, 1, 7, -21, 16, 0, 19, 7, 36, 26, 33, 9, -9, 13, -3, 18, -7, -8, 15, -17, 61, 73, 30, 47, 45, 81, 55, 57, 59, 13, -7, -26, -17, 26, 35, 31, 47, 32, 34, 63, 0, -17, 11, 9, -7, 17, -5, -6, 60, 53, 61, 51, 65, 28, 6, 52, 38, -14, -18, -16, 8, 13, 26, 22, 11, 7, 22, 12, 1, 6, 17, 4, 16, 12, -13, 0, 47, 39, 61, 42, -8, -20, -38, -18, -12, -20, -10, 14, 20, 34, -10, 9, 16, -13, 35, 8, 15, -42, 2, -11, 0, 15, 10, -30, 25, 16, -15, -25, -57, -42, -37, -29, -32, 1, 19, 24, 11, 5, -16, -5, -26, -50, -12, 4, -5, -24, 17, -7, 3, -14, 19, -65, -13, -28, -45, -85, -45, -22, 14, 5, 8, 39, 2, -8, -16, -16, -26, -25, -61, -63, -10, 20, 26, -22, -15, -15, 0, 15, -3, -11, 35, -37, -28, -20, -32, 15, 13, 25, 16, 31, 42, 7, -9, 0, -34, -16, -9, -2, -16, 5, 24, 14, 2, -9, 17, 12, 23, -31, 11, -19, -37, -30, -42, -9, 0, -6, -2, -13, 11, -4, -12, -36, -15, -36, -13, -6, -26, 6, -17, -12, -1, -13, -13, -19, 50, 0, 3, -4, -37, -54, -49, -40, -43, -23, -14, -16, 12, 10, 1, 25, 26, 13, 11, 16, -39, -31, 5, 29, 5, 17, 14, 7, -2, -10, 12, 6, -17, -47, -26, -24, -14, 5, 16, 20, 15, 26, 49, 71, 48, 43, -7, 12, -12, -5, 32, 39, -5, 7, -16, 5, -37, 57, 51, 54, -3, 7, 18, 22, 25, 30, 74, 46, 48, 55, 35, 54, 60, 71, 23, -29, -7, 8, 15, -4, -8, -15, 7, -4, 14, 48, 87, 65, 67, 38, 55, 65, 67, 49, 44, 37, 39, 55, 78, 40, 19, 36, -6, -16, 11, -3, -18, -52, -13, -18, 20, -20, 37, 54, 94, 84, 57, 49, 75, 69, 84, 60, 4, 28, -15, 9, 40, 8, -2, -11, -8, -26, -19, -12, -3, -45, -9, 9, -14, -4, 45, 75, 83, 73, 67, 104, 102, 58, 67, 16, 46, 10, -11, 8, 19, 5, -26, -3, -31, -25, -19, 7, 33, -41, 12, -1, 17, -14, 37, 16, 94, 62, 34, 46, 82, 97, 72, 18, 22, -9, -24, 22, 22, 2, -5, 7, 16, -9, -17, 26, 16, -33, 6, -4, -20, -14, -3, 46, 56, 48, 11, 32, 64, 43, 22, -15, -12, -32, 7, 9, 43, -6, 11, 32, 22, 38, 63, 39, 48, -10, -1, -17, -18, -3, -10, 27, 24, 32, -1, 8, 10, 32, 8, 3, -3, -2, -18, 52, 17, 11, 19, 36, 33, 4, 73, 47, 19, 26, -4, -7, -6, 2, -6, -7, 8, -23, -20, -22, -24, 23, 19, -10, -16, 16, 35, 24, 25, -10, 35, 48, -1, 23, 70, 53, 94, -15, 8, -7, -8, -19, -26, 33, 6, -6, -9, -5, 3, 42, 35, -8, -13, 18, 10, 7, 19, 0, 15, 40, 47, 48, 58, 34, 67, -7, -8, 11, -20, -15, 30, 23, 57, 0, 21, 18, 29, 5, -31, -23, -24, 18, 14, -11, 5, 12, -3, 6, 23, 45, 26, 6, -4, -2, -18, -12, 9, -12, -9, 59, 47, 45, 22, 15, 27, 28, -26, -44, -36, -22, -28, -24, 27, -8, -1, 21, 45, 50, 49, 30, 3, -1, 1, -14, 5, 15, -10, 66, 73, 63, 69, 49, 32, 18, 13, 14, -29, -41, -11, 10, 0, 9, -6, 2, 55, 33, 30, 27, 27, 2),
  79 => (13, 11, -17, -14, 19, 11, 4, 8, -5, -2, 13, 20, -7, -5, -13, 0, 25, -14, -19, 13, -39, -31, -21, 20, 18, 1, 16, -15, -1, -5, 19, 9, 14, -13, 8, -3, -9, -8, 6, 8, 13, 47, 44, 36, 44, -2, 5, -12, -24, -18, -22, 43, 33, 0, -4, 11, 7, 18, -5, -16, 20, -7, -10, -14, 4, 19, 4, 22, 73, 48, 55, 33, 8, -17, -27, -26, -72, -8, 16, 48, 5, -33, 12, 13, -1, -20, 17, -10, -13, 15, -2, 7, 2, 14, 36, 41, 49, 49, -23, -40, -20, -69, -49, -21, -25, -25, -5, -15, -11, 24, -10, 20, -12, -5, 17, -1, 9, -2, 17, -16, 6, 17, 24, 33, -16, -14, -39, -41, -61, -47, -12, 2, 0, -21, -20, 18, -13, -1, 17, -5, 6, -1, 2, 15, -4, -5, 14, -14, 10, 30, 19, -31, -27, -14, -23, -12, -23, -11, -13, -15, -12, -27, 11, 26, 62, -21, 5, 15, 21, -14, -19, 9, -21, 10, 17, -18, 14, -1, -20, 7, 17, 51, 25, -9, -36, -38, -42, 4, -9, -13, 0, 14, 46, 31, -24, 8, 12, -16, 4, -15, 11, 15, 0, -7, -27, 4, 57, 40, 38, 53, 8, -7, -34, -6, -15, 14, 7, -17, -13, 33, 18, 17, -24, 8, -13, 10, 20, 12, -15, -6, -15, -10, -31, 22, 35, -3, 9, 10, 37, 1, -39, -23, -6, 4, 4, 16, 44, 44, -10, 16, 11, -7, -7, -12, -13, -2, 13, 1, 6, -12, -41, 2, -3, -42, -23, 12, -26, -47, -36, -37, 9, -1, 1, -6, 35, 18, 9, -14, 5, -4, -2, 18, 17, -2, 4, -11, -21, 12, -45, 6, 16, -30, -19, -7, -18, -33, -32, -2, 20, -9, -27, 1, 26, 18, 4, -24, -7, -2, -7, -11, 8, -2, 13, -16, 1, -21, -71, -65, -4, -18, -11, -25, -43, -92, -48, 7, 16, 2, 14, 38, 27, -3, -18, -49, 13, -17, -8, 14, -11, 15, -11, -9, 0, -14, -67, -86, -78, -35, -57, -89, -119, -106, -23, 46, 30, 17, -4, 22, 6, -6, -24, -50, 8, 12, 7, -4, -1, -15, 10, -1, 14, 7, -55, -98, -77, -72, -76, -102, -87, -49, -7, 59, 15, 26, 18, -4, -10, 19, 17, -4, -8, -7, -14, -11, 19, 19, 6, 5, 16, 0, -23, -58, -63, -79, -74, -66, -58, -20, 35, 45, 57, 44, 17, 19, 11, 14, 11, 7, -19, -5, -14, 16, 3, 1, -22, -20, -6, 25, -38, -40, -62, -124, -59, -42, 13, 31, 44, 47, 36, 23, 47, 26, 12, -12, -32, 17, 5, 27, 12, 8, 1, -3, -2, -31, -6, -25, -5, -29, -41, -38, -27, -12, 13, 36, 27, 19, 31, 9, 12, 5, 15, -29, -35, -10, -3, 4, 1, 3, 16, 17, -7, 1, 7, -26, 3, -29, -33, -30, -13, 8, 41, 33, 17, 30, 19, 42, 10, 31, 15, -9, -30, -15, -9, -10, 15, -13, -20, 2, -15, -11, -3, 10, -9, -31, -51, -8, 3, 7, 24, 28, 43, 38, 32, 23, 32, 35, 33, 18, 18, -7, -23, -11, 10, 16, -7, -4, 2, 7, -25, 5, -29, -41, -58, -36, -15, -10, 1, 26, 28, 0, 46, 21, 3, 13, 16, 1, 6, -18, 12, 20, 7, 14, -9, -11, -18, 7, -32, -44, -51, -96, -54, -59, -1, 9, 17, 56, 35, 24, 24, -4, 21, 0, 18, -11, -9, -25, -52, 14, -14, -8, -6, 14, 14, -16, -46, -85, -47, -83, -53, -12, 5, 32, 48, 56, 39, 3, 23, 10, 11, 26, 21, -20, -23, -29, -38, 0, -17, 4, -16, -12, -19, -8, -35, -65, -73, -54, -24, -31, 8, 39, 7, 45, 28, 5, 15, 9, 34, 24, -13, -11, -15, -45, -31, 31, -16, -5, 0, 6, -9, -3, 0, -17, -6, -38, -29, 6, 46, 64, 24, 27, 18, 4, 7, 35, 23, -1, 0, -16, -11, -46, -29, -9, 1, -15, 7, 7, 15, 26, -7, 1, 22, 12, 34, 71, 80, 77, 55, 31, 21, 8, 25, 30, 11, 28, -13, -2, -37, -43, -7, 16, -17, -3, 3, -19, 14, -10, -4, -34, 23, 10, 36, 15, 58, 52, 28, 37, 5, -14, -15, -5, -2, 0, 9, -28, -55, -55, -36, 20, -9, 4, 17, 10, -16, 11, 16, 6, 15, 5, 9, 9, 27, 36, 29, 22, 29, 17, 3, -10, -50, -23, -9, 15, -8, -26, 1, 31, 7, 17, 8, -7, -17, 11, 22, -4, -14, -17, -9, 30, 39, 43, 18, 35, 28, 27, -10, 25, -7, -4, -19, 21, 27, 17, 14, 14),
  80 => (3, 0, -15, 20, 12, -5, -1, 10, -3, -15, -17, 11, -15, 6, 2, -35, -1, 14, 15, -35, -38, -14, -12, -14, 6, 1, -1, 9, 17, 7, -6, -11, 11, -1, -15, 19, -4, -9, 12, -19, -31, -2, -12, -29, -4, -2, -14, -22, -14, -23, 34, 57, 29, 19, -20, -18, -5, -3, -12, 12, 6, -5, 19, 4, 6, 4, 10, -28, -17, -41, -41, -33, -2, -27, -10, -23, 12, 39, 42, 49, 24, -5, 2, 10, 15, -17, 19, -18, -5, -2, 8, 6, -12, -15, -8, 10, 8, 6, 15, -27, -18, -25, -20, 20, 19, 31, 49, 38, 35, 18, -6, 3, -17, -11, -16, -12, 13, -8, -1, -10, 0, -6, -13, 14, -5, -18, -10, -30, -27, -22, -17, -32, -31, 18, 35, 42, 26, 58, -19, 19, -10, 21, -19, -15, -21, -16, -14, 11, 21, -8, -4, 21, -42, -44, -25, -21, 7, -30, -66, -52, -16, 21, 27, 57, 34, 62, 13, 11, 11, -17, 9, 4, 2, -18, -14, 16, 20, 9, -36, -21, -55, -42, -28, 13, -11, -28, -27, -13, 3, 14, 25, 33, 33, 13, 18, -18, 15, 4, 13, -6, 14, -8, 24, 36, -18, -19, -54, -44, -67, -59, -25, -27, -29, -34, -52, -27, -19, -28, 14, 35, 3, -8, 24, 22, -6, -19, -4, 9, 11, 11, 23, 8, -14, -62, -68, -27, -44, -26, -40, -28, -31, -29, -35, 11, -22, 15, -2, 7, 5, 34, 4, 21, -5, 2, 0, -7, 21, -10, 45, 27, -69, -77, -71, -28, -14, -13, -28, -32, -40, -65, -69, 17, 0, 6, 21, 24, 5, 25, 15, -3, 15, -15, 7, 1, 14, 5, -12, -3, -51, -27, -1, -26, -17, -34, -29, -38, -43, -72, -95, -22, -34, 9, 41, 29, 4, 29, -27, 14, -10, 6, 13, -13, -15, -11, 8, -36, -23, -31, -4, 7, -1, -38, -16, -20, -22, -30, -36, -53, 5, 21, -8, 29, 2, -1, -19, 24, 11, 16, 11, -16, -16, -7, -29, -22, -39, -17, 18, 3, 18, 2, -2, -60, -30, 6, -36, -37, 20, 46, 14, 8, 21, 12, 10, 22, 21, -4, -13, 7, 17, -4, 0, -25, 0, -4, -22, 24, -9, -9, -25, -50, -83, -26, -8, 13, 36, 45, 17, 30, 30, 22, -7, 43, 15, -18, -1, -13, -31, -20, -19, 9, 15, 6, -15, 31, -18, -24, -21, -49, -47, 20, 60, 58, 70, 69, 32, 18, -13, -11, -26, 42, 2, -13, -15, -15, 9, 3, 36, 38, 34, -23, -43, 18, 4, -23, -10, -33, -20, 67, 67, 40, 54, 56, 10, 32, -27, -36, -25, -15, 18, 0, -13, -14, -9, 43, 31, 52, 36, -7, -22, -3, 14, 7, -13, -44, -17, 11, 55, 30, 40, 26, 20, -17, -4, 1, 0, 8, -4, -9, 20, -12, 14, 24, 40, 67, 30, 20, -5, 0, 26, 12, -7, -17, -13, -18, -2, 22, 43, 41, 9, -27, 1, -14, -19, 0, 21, -6, -20, -13, 29, 56, 52, 18, 36, 41, 39, 49, 9, 1, -38, -42, -55, -18, -6, 7, 29, 33, 13, -27, -15, -30, -10, -9, -9, 0, -19, -3, 11, 39, 21, 24, 26, 1, 33, 17, 13, 12, -36, -31, -42, -20, -8, 23, 19, 27, -20, -57, 5, -10, -20, 20, -11, 11, -7, -1, 27, 29, 65, -8, 10, 20, 24, 9, 15, 18, -40, -22, -64, -40, -23, -12, -2, -2, 10, -15, 19, 10, -36, 4, -7, 10, -15, -16, 4, 42, -5, -54, -32, -61, -15, 45, 12, 18, -16, -25, -35, -46, 15, 15, -11, 3, 23, -14, -4, -8, -46, -38, 4, 19, 4, 20, 12, 32, -14, -49, -51, -60, -30, 24, 5, 11, -41, -25, -31, -1, -13, 27, 10, 17, 6, 9, -18, 15, -77, -35, -5, -21, -8, 11, 25, 41, 6, -45, -56, -48, -12, 3, -11, -5, 34, -12, 14, 17, 37, 31, -11, 17, 16, 20, 13, -13, -50, -9, 0, -1, 14, -19, 2, 50, 21, -45, -50, -47, -22, 27, 16, 3, 11, 30, 32, 28, 18, 28, 2, 23, 2, -30, -19, -7, -13, 13, 7, -1, 0, 8, -16, 3, -18, -51, -79, -66, -19, -10, 59, 43, 13, 17, 31, -3, 27, 7, 25, 16, 18, -22, -31, -33, -64, 7, 7, -6, -17, 11, 0, 11, 1, -3, -38, -49, -19, -10, 29, 47, 8, -1, 26, 30, 44, 6, 48, 32, 18, 19, -14, -37, -33, -1, -9, -15, -9, -1, -1, 23, 14, -15, -36, -30, -31, -13, -12, -32, 0, -10, 8, 2, -23, 28, -18, 7, 9, 1, 28, -4, 12, 6),
  81 => (19, 20, -16, -9, -5, 19, 3, 1, 10, -12, 18, -9, -15, 10, 18, -1, -22, -8, 17, -42, -34, -38, 1, 15, -12, -10, 17, -20, 16, -7, 16, 16, 1, -4, 7, 9, -7, 6, 20, -18, -34, -25, -4, 3, -25, 8, -5, 0, -12, -39, 9, -12, -8, -5, 11, 0, -13, 20, -5, -7, 19, 4, -9, 8, 14, -46, -32, -2, -2, -36, -21, -4, -8, 26, -11, 33, 7, 1, -56, -38, -53, 9, -16, 19, 3, -5, -11, 5, 8, -2, -20, -1, -23, -14, -8, 1, -4, 10, 2, 12, -24, -6, -20, -51, -26, -23, 29, -23, -1, -24, -1, 3, -9, -1, -11, 1, -13, 18, -9, 10, -12, -19, -37, -90, -57, 13, 48, 18, 11, -23, -68, -52, -34, -32, -9, -2, -10, -10, -9, 9, -16, -9, -20, -10, -17, 11, 0, -12, -25, -52, -99, -112, -63, 16, 12, 14, -41, 9, -51, -94, -25, -35, -10, -18, 1, -7, 8, -2, -3, 13, -20, 5, -1, -19, 12, -10, -27, -75, -85, -87, -52, -1, -13, -17, -7, -24, -24, -50, -14, -22, 21, -14, 11, 50, 9, 16, 2, 7, 5, -15, 1, -20, -6, -41, -37, -71, -78, -59, -45, -14, -31, 22, -40, -25, -46, -1, 19, -5, -28, -20, 30, 24, 40, 9, 10, 5, -1, -7, 2, 20, -13, -15, -66, -56, -64, -44, -22, -48, -64, -16, -30, 7, -13, 46, 30, 40, 20, 3, 52, 87, 50, 60, 3, 14, -7, -6, 3, -17, 26, -65, -81, -48, -50, -41, -21, 7, 16, 47, 9, 6, -3, 27, 12, 19, -4, -4, 21, 47, 74, 59, 14, 11, 1, 20, 8, 48, 5, -44, -11, 6, 33, 17, 64, 89, 54, 60, 12, 23, -8, 17, 26, -7, 13, -23, 16, 33, 62, 44, -15, -15, -9, -18, 7, 55, 6, 34, 67, 98, 62, 24, 82, 63, 15, 21, 37, 35, 28, -2, 37, 29, 28, 61, 39, 36, 25, 9, -1, -10, 11, -7, 38, 32, -2, 4, 49, 20, 35, 44, 53, 86, 22, 36, 14, -14, 3, -1, 4, -8, 27, 57, 23, 0, -7, 37, -3, -3, -6, 6, 4, 19, 6, 36, -5, 25, 38, -8, 58, 49, 24, 0, -4, 3, 26, 6, -10, 28, 14, 30, -7, -44, -7, 26, -16, 6, -6, 19, -6, 8, -5, 10, 3, -13, 15, 8, 34, 39, 17, 29, 26, 46, 46, -20, -1, 20, -16, -2, -14, -6, -25, -10, 3, -9, 16, -8, 5, 12, -22, -8, 18, 28, 13, 38, 37, 5, 12, 6, -1, 18, 30, -1, 25, 16, -12, -16, 4, -9, -42, -8, 5, 7, -20, -10, 43, 17, -2, 53, 26, 9, 33, 37, 26, 9, 17, 27, -28, -23, -8, -13, 22, 13, -14, -47, 6, -7, -11, -12, -3, 2, 3, -1, 14, 21, 44, 35, 13, -1, 21, -18, -34, -13, -28, -29, -69, -31, -2, -27, -49, -20, -31, -40, -12, -23, -38, 9, -18, -16, -15, 19, 43, 22, 41, 30, -4, -2, 16, -33, -46, -11, -7, -52, -59, -25, -44, -62, -65, -46, -58, -61, -3, 7, -33, 33, -12, 20, 1, 2, 36, 2, 51, 23, 34, -9, 24, -3, -58, -1, -18, -21, 16, -49, -57, -29, -47, -39, -58, -64, -32, -10, -19, 35, -15, -14, -11, 5, -32, -31, -34, -9, 22, -4, 14, -34, -39, -33, -51, -2, 21, -32, -60, -41, -38, -46, -48, -37, 4, 8, 13, 1, 15, -16, 11, -19, 8, -22, -71, -36, -9, 2, 28, -16, -33, -2, -5, -3, 12, 1, -15, -9, -6, -35, 10, 6, 10, -17, -8, 17, 13, -17, -12, 0, -19, -25, -42, -20, -34, 8, -3, 14, 6, 23, -5, 1, -11, 36, -15, 40, 14, -15, -28, -13, -13, -17, -40, 11, 6, 20, -15, 0, -22, -25, -1, 34, -16, -9, -13, 21, 17, 9, -29, -39, -31, -35, -53, -38, 11, 11, -7, 5, -7, -3, 25, -5, 2, 2, 4, -17, -19, -15, 10, 11, 41, 17, -34, -39, -15, -18, -53, -50, -90, -27, -62, -55, -38, 4, 20, 33, -23, -17, 12, 25, 5, -6, 6, 11, -13, 38, 18, 38, 22, -10, -35, -47, -8, 3, -19, -16, -17, -55, -37, -4, 7, 14, -10, 13, 3, -25, -1, 16, -3, 3, -10, -1, 9, -42, 7, 22, 52, 29, -1, -35, -21, 9, -8, 8, 13, -6, -10, -6, 47, 30, 18, -21, 27, -4, -42, 32, -5, -11, -13, 8, -18, -15, -28, -63, -58, -10, 0, -36, -58, -100, -25, 9, 17, -3, -5, 19, 18, 10, 10, 6, 15, 0, 6, 16),
  82 => (15, 1, 11, 2, 3, -14, -6, 19, 2, -4, 19, -12, 3, 12, 15, -10, -54, -22, 9, 10, -6, -2, -14, 11, -5, -12, 7, 6, -1, -1, 6, 16, -10, 3, -10, -16, 18, -19, 8, -16, -19, -29, -22, 7, -12, -12, 4, 10, -10, -11, -19, -18, -5, -13, -18, -14, 15, 4, 5, -2, -17, -13, 4, -2, 16, -22, -7, -20, 2, 7, 24, -1, -18, -37, -29, -37, -36, -18, -14, -11, -32, -16, -5, 1, 10, -20, 9, -7, -6, 7, -9, -12, 10, -20, 20, -16, -18, -12, -28, -37, -44, -46, -44, -44, -56, -35, -9, -36, -15, -1, 15, -6, 16, 3, 14, 19, -19, 5, 10, 1, -25, 3, -13, 10, 2, -24, -9, 3, -4, -55, -13, -27, -43, -15, -22, -17, -12, 24, 9, -11, 9, -8, 9, 10, 4, -1, 11, 8, 36, 19, 4, 11, -17, 1, -28, 21, -20, -10, -13, -27, -7, -8, -14, 14, -6, -4, 2, -3, 4, 17, 16, -4, -10, -12, -26, -37, 12, 48, 1, -15, 11, -23, -17, -26, -7, -21, -3, -34, -8, -21, 8, 8, 7, 19, 1, 14, -6, -14, -3, 10, -16, 3, 2, -59, -18, 2, -16, -5, -4, -33, -28, -20, 2, -13, 12, 19, 5, -11, 12, 17, -10, 5, 8, -6, 13, 0, -13, -17, 14, -21, -18, -32, -23, -20, -19, 8, 10, 4, 3, 10, -23, -14, 27, -10, -4, -9, 4, 11, -20, 2, 27, 53, 2, -17, -3, -19, -20, 8, -5, -30, -35, -3, -2, -17, 16, 11, -39, -46, -3, 11, 44, 9, 20, -5, -23, -22, 39, 14, 31, 74, -16, 1, -16, -21, -2, 5, -7, -17, 3, -19, 0, -30, -7, 4, -4, 6, 38, 25, 43, 44, 33, 11, 8, 25, 14, 13, 6, 35, 19, -11, 20, -10, 1, 18, -20, 12, 30, 50, 19, 22, 14, 13, 8, 20, 19, -7, 15, 34, 33, 25, 4, -25, -3, 4, -17, 17, -11, 20, 9, -7, 15, 26, 51, 60, 55, 63, 23, 12, 27, 23, 38, 5, 22, 0, 0, 23, 26, -13, 21, 14, -13, -15, 14, -11, 11, 19, -13, -14, 21, 36, 41, 57, 68, 65, 47, 50, 31, 52, 20, 19, -19, -45, -3, 3, 8, -6, -38, 14, 15, 5, -19, -1, 1, 14, 11, -12, -30, 19, 68, 9, 25, 36, 0, 2, -7, -17, -27, -45, -32, -55, -15, -17, -33, -16, -6, 8, 5, 37, -11, -42, 12, 14, -6, 14, 11, 7, -2, 0, -29, -53, -67, -50, -75, -16, -41, -5, -4, -41, 2, 10, -7, 2, 16, 16, 18, 37, 4, -22, -15, 6, -9, 12, 16, 2, -63, -52, -25, -75, -4, -1, 12, 25, -7, -3, -6, -33, -32, 23, 23, -14, -11, -7, -3, 32, 47, 30, 1, 19, 1, 4, -9, -17, -80, -30, -41, -55, -43, -17, 4, 11, -4, -30, -30, -36, -64, -29, -46, -9, -10, 16, -6, -25, 17, 1, 20, -15, 8, -16, -3, -26, -15, 12, -30, -67, -65, -57, -72, -32, -15, -43, -39, -53, -45, -49, -14, -4, -29, -21, 18, 2, 10, -13, 0, -16, -3, -10, -1, -18, -29, 15, -2, -56, -55, -78, -85, -85, -81, -46, -65, -68, -65, -22, -33, 26, 39, 9, -22, -7, -1, -27, 3, -11, -15, -14, -41, -43, -29, -18, 16, -39, -27, -31, -69, -127, -87, -50, -66, -53, -41, -31, -7, -10, 21, 27, -10, 11, -9, 8, 19, -4, -17, -2, -9, -35, -13, 24, 26, -4, -12, -14, -2, -28, -18, 8, -22, 3, 12, 14, 45, 0, -18, 20, 56, 47, 36, -4, 14, -16, 18, -6, 24, 18, 2, -4, 41, 21, -16, -5, -3, 14, 39, 38, 45, 46, 28, 54, 22, -28, 10, 13, 25, 50, 34, 40, 16, 16, -13, 2, 14, 30, -13, 28, 24, 20, 28, 17, 13, 53, 28, 45, 38, 70, 56, 44, 20, -7, 16, 38, 41, 30, 23, 9, -4, 7, -3, -12, 10, 28, 14, 1, 46, 48, 27, 29, 56, 41, 23, 2, 20, 52, 52, 58, 24, -12, -1, 1, -13, 14, 18, 17, -9, -12, -21, -11, 12, 41, 16, 20, 35, 9, 40, 36, 33, 58, 32, 20, 32, 58, 28, 29, 40, -4, 14, 13, 10, -31, 1, 19, 17, 1, 11, 7, 35, 20, 44, 50, 67, 13, -17, 4, -3, -11, -1, 22, 51, 74, 29, 62, 17, 22, -17, 4, -26, -16, 30, 5, 11, 0, -9, -19, -17, 3, 12, -3, 9, 27, 27, 9, 13, 10, 30, 21, 39, 45, 37, 13, 5, 10, 0, -16, -29, -10, 25, 56),
  83 => (-15, -4, -13, 16, -18, 3, -5, -4, 14, 15, 10, 17, 6, 17, 41, -17, 47, 33, 33, 40, 19, -10, 5, 14, 5, -18, 18, -3, 19, -20, -2, -17, -20, 20, -5, 19, -13, -16, -37, -12, 26, 51, 16, 22, 42, -4, 43, -18, -4, 17, 10, 12, -13, -17, 17, -4, -3, -12, -2, 2, -4, -12, -13, 16, -7, -7, 32, 52, 6, 38, 31, 39, -58, -98, -21, -35, -43, 10, 23, -12, 5, -5, 1, 12, 6, -19, 12, 17, 18, -10, -16, -3, 29, 22, 41, 34, 25, 8, -34, -35, -101, -109, -78, -23, -12, -32, 8, 6, 8, 7, -10, 20, 0, 17, -20, -4, -13, 4, -7, -27, -7, -39, -11, 25, 57, 28, -1, 2, -42, -112, -135, -58, 1, -53, -2, 6, -4, -11, 14, 11, 8, 19, 3, 14, -8, -19, 2, 28, -27, 13, 41, 55, 46, 21, -28, -23, -37, -51, -111, -68, -55, -61, 0, 16, 19, -11, 17, 10, -7, -5, -13, -3, 11, 9, -17, 36, -19, 10, 28, 17, 33, 48, -1, -5, 18, -68, -155, -141, -95, -80, -11, -1, -19, 13, -5, -21, -19, -1, 8, 19, -6, -11, 11, -23, -14, 12, 5, 44, 65, 29, 50, 29, 11, -5, -85, -128, -119, -54, -41, -8, -14, 18, 5, -15, -20, -11, -1, 3, -13, -11, 13, -8, -39, -8, -47, -1, 21, 20, 66, 32, 46, 8, -34, -85, -106, -80, -97, -60, -14, -21, 10, 14, 17, 6, 11, 3, 6, -9, -22, -60, -23, -46, -42, -21, -5, 15, 48, 55, 21, 3, 5, -6, -67, -88, -69, -68, -9, -21, -16, -17, -5, 0, 4, 16, -7, -29, -42, -62, -51, -52, -1, -22, 8, 7, 5, 44, 2, 6, 3, -21, -39, -62, -70, -77, -27, -24, -27, 7, -10, -9, -2, 16, 1, -35, -38, -38, -20, -15, -4, -4, 24, -13, 0, 51, 6, 20, 23, -23, -12, -5, -31, -54, -47, 1, 6, -3, 12, 6, -20, -19, 20, -26, 29, -11, 2, -15, -5, -12, -3, 11, 24, 53, 18, 29, 9, 11, 20, 26, 13, -26, -48, -46, -25, -1, 17, -3, 8, -10, -8, -19, 72, 24, 7, -32, -39, 6, -3, 2, 13, 28, 53, 41, 9, 47, 37, 52, 9, -14, -1, -2, -21, -1, 1, -17, -14, -7, 47, 27, 37, 11, -2, 6, -30, -24, -25, 30, 3, 3, 43, 28, 16, 39, 39, 5, 12, -4, 14, -13, -12, 2, 20, -9, -7, -8, 17, 63, 8, 15, -11, -17, -32, -21, -13, 5, 4, -37, 4, 7, 13, 27, -8, 6, -38, -14, -21, -16, -24, -30, 14, -1, -9, -9, 28, 4, 7, -7, -30, -42, -49, -39, -36, -13, -6, -38, -57, -36, -10, -20, -30, -1, -37, -51, -31, -20, -22, -15, 8, -17, 12, -5, 8, 7, -11, -52, -39, -51, -44, -30, -27, -4, -17, -16, -29, -24, -73, -21, -37, -38, -13, -37, -39, -22, -49, -7, -3, -18, 13, -17, -4, 33, -17, -2, 19, -6, -2, -20, -30, -5, 7, -39, -25, -42, -51, -12, -31, -18, -39, -49, -33, -51, -49, -13, -14, -7, -20, -4, -19, 36, 6, 4, -4, 20, 12, 11, -44, 9, 21, 9, 4, -1, -22, 0, -33, -22, -34, -25, -65, -59, -15, -5, 15, -5, 5, 7, 16, 23, 26, 53, 30, 26, 60, 45, 23, 74, 34, -10, 24, 29, 4, -15, -3, 27, -10, -10, -55, -42, -36, 11, -19, -16, -18, 8, 9, 34, 56, 46, 15, 14, 39, 19, 21, 41, 26, 11, 23, -10, 7, 18, 39, 30, 34, -18, -19, 2, 0, -12, 14, 7, 1, 0, 14, 8, 9, 18, 13, 26, 37, 11, 14, 48, 9, 40, 34, 28, 10, 6, 35, 45, 50, 25, -13, 30, 7, 14, 17, -3, -14, -13, 69, 42, 24, 14, 37, 10, 19, 32, 28, 36, -13, 15, 24, 17, 1, 1, 20, 13, -4, -11, -18, 16, 12, 22, -17, -3, 9, -4, 59, 60, -7, 21, 47, 24, 5, 27, 35, 25, 10, 8, -10, 10, -8, -15, 20, 27, 1, -2, -5, -13, 13, 25, -12, -17, -12, 8, 26, -13, -29, -37, -11, 7, -3, -19, 14, 7, 18, -8, -39, -31, 12, 14, 4, 11, 13, 17, -2, -3, -6, 43, -8, -12, -15, 7, 9, -5, 13, 11, -32, -28, -40, -32, -34, -78, -43, -22, -10, -37, -20, -29, 2, 13, 27, 22, 29, 15, -2, 48, -13, 3, -1, -16, 17, -3, -32, -37, -40, -31, -26, -40, -35, -28, -23, -9, 0, 2, -11, -25, -30, 14, 32, 30, 42, 56, 69, 30),
  84 => (6, 6, 0, 2, 5, -6, -5, -5, -4, -17, -6, 19, -11, -12, 8, -30, -72, -51, -26, -16, 3, 5, -9, 14, 2, -1, -7, 19, -6, 16, 2, -14, 11, 4, 17, 11, -7, -18, 24, 67, 41, 30, 30, -7, 39, 33, 11, 36, 7, 10, 56, -28, -38, 5, -9, -19, 10, -8, -13, -7, -8, -5, -18, -18, -10, 58, 26, 70, 41, 32, 84, 57, 49, 55, 41, 31, -1, -17, -40, -8, -45, -41, -10, 2, -4, 8, 12, 12, 2, -19, 2, -3, 38, 33, 56, 46, 5, 51, 48, 5, 19, 3, 6, -30, -28, 11, -19, -29, -14, -25, -11, 0, -3, 15, -13, 13, -20, 0, -20, 27, 42, -8, -24, -15, 4, -22, 15, -5, 38, 25, 4, -6, -13, 26, 61, 47, 0, -12, 5, -12, -4, 12, -15, 15, 20, -6, 1, 28, 2, -22, -30, -1, 3, 24, 28, 37, 14, 10, 3, -9, 1, -1, 45, 21, -3, -5, -7, 1, -9, -13, -16, -7, 7, -1, 36, 57, -7, 36, 37, 66, 39, 28, 45, 14, 9, 11, -17, 10, 26, 23, 68, 39, 45, 10, -14, 18, 6, 5, -5, -11, 1, 8, 53, 41, 23, 67, 38, 15, -18, 2, 25, 9, 9, 6, -8, 16, 6, 27, 24, -8, 28, 14, -1, -8, 8, 9, -18, -16, -3, -16, 21, 31, 46, 38, -44, -28, -38, 1, 28, 42, 5, 1, 28, 19, -9, 3, 9, -17, 33, 14, -23, 4, -12, 2, 7, 12, -18, -19, -26, 20, 12, -15, -50, -13, -18, -15, 0, 21, 10, 9, 8, 34, 34, 36, 2, -21, -19, 4, 47, 70, 7, 10, -3, 0, 5, -10, 9, 14, 18, -22, -5, 28, -28, 16, -11, -14, -3, -23, -45, -52, -13, -29, 11, 12, -57, -12, 29, -3, 6, -8, 20, 8, -10, -30, 19, 11, -12, 1, -22, 2, 17, 7, 15, 23, 1, -17, -31, 1, -25, 9, 2, 5, -11, -66, 14, -46, -21, 4, 3, 9, 21, 39, 56, -13, -16, -20, -34, 17, 13, 9, 1, -10, -8, 1, 16, 10, 8, -15, 8, 4, -9, -29, -13, -37, 4, -15, 18, 0, 51, 20, 19, -22, -16, -12, -23, 10, 9, -4, 9, -5, 18, 30, -9, 18, 31, 11, 10, 24, -34, -16, 9, 4, -13, 1, -10, 20, 5, 15, 14, 13, -15, 11, 6, -11, 1, 23, 48, 13, 51, 79, 40, 58, 33, 31, 2, -1, -11, -36, -28, 38, -19, 4, -9, 7, -8, 30, 6, 17, 35, 66, 47, 26, 65, 64, 35, 63, 77, 77, 41, 87, 67, 7, -14, 1, 3, -40, -6, 57, 3, -5, -1, 11, 28, 29, 26, 67, 65, 77, 83, 82, 89, 69, 67, 98, 76, 58, 41, 45, 35, 29, 13, 25, -24, -35, 12, 29, 16, 11, -15, 10, 12, 21, 74, 69, 106, 88, 101, 91, 82, 86, 79, 52, 63, 18, 2, 6, 11, -13, -15, 10, 3, 19, 20, 18, 9, -17, -4, -13, 24, 51, 62, 64, 61, 42, 56, 24, 28, 26, 8, 40, -13, 7, -5, -8, 3, -17, -9, -17, 5, 19, 20, -4, 17, 10, 10, 13, 16, 39, 58, 26, 24, 42, 25, 28, -11, -12, 13, -20, -24, 14, 2, -12, 8, 13, 14, -3, -25, 16, 12, 30, 9, -11, -16, 5, -22, -20, 23, -9, 16, -13, 28, -1, -2, -18, -29, -35, -13, 5, -8, -11, 1, -6, 42, 64, 34, 35, 34, 43, 7, 8, -8, 1, 9, 1, 21, 2, -21, -9, 39, 15, 5, 22, 7, -14, 0, -3, -12, -17, 6, 18, 33, 85, 88, 34, 60, 29, -19, -4, -4, 15, 37, -21, -15, 4, 5, -19, 30, 43, 46, 23, 15, -10, -9, 14, 4, -1, 28, 58, 37, 85, 52, 67, 15, -29, -18, 14, -20, -4, 36, 2, 40, 26, -14, 12, -4, 22, 36, 40, 28, 29, 42, 28, 27, 50, 73, 64, 42, 46, 31, 24, 44, -34, 19, 11, -4, -11, -18, 5, 50, 14, 23, 23, 25, 49, 62, 66, 55, 57, 33, 38, 67, 67, 72, 69, 53, 12, 21, 7, 16, 4, -13, -11, 18, -9, -10, 57, 32, 4, 9, 4, 10, 48, 42, 20, 5, 24, 31, 11, 34, 73, 50, 65, -2, 25, 20, -27, 7, -19, 19, -2, -16, -16, 1, 52, 70, 25, 14, -5, 6, 33, 22, 18, 46, 4, -3, -10, 9, 0, -1, -1, -9, 21, 4, -41, -25, -50, 10, -18, -17, -3, 0, 5, 27, 71, 31, 25, -11, 1, 21, -10, 13, 61, 11, -5, 2, 7, -21, -47, -65, -38, -34, -29, -20, -17),
  85 => (18, -14, -1, -19, 20, 16, -1, -17, 9, 5, -3, -8, 16, -13, -19, 10, 21, 58, 24, 59, 42, 5, -19, 18, -2, -20, -14, 17, 4, -3, 1, 14, 1, -20, -12, -19, -21, -12, -4, 15, 11, -50, -20, 25, 2, 38, 57, 79, 57, 61, 17, -11, -5, 3, 7, 6, 16, -15, 12, 17, -14, 20, 8, 3, 8, -20, -3, -23, -56, -5, -21, 13, 28, 54, 61, 35, 48, 31, -28, 16, -24, -6, -3, 6, 10, 18, -7, 3, -3, 6, 9, -17, -7, 11, -10, 2, 18, 44, 44, 34, 19, 46, 57, 39, 17, -20, 38, 0, -64, -33, 18, 7, -19, 4, 14, -17, -19, 19, -5, 7, 14, -32, -5, -16, 45, 52, 59, 31, 18, 27, 84, 56, 8, -22, 36, 21, -32, -13, -14, 11, 11, -1, -21, -10, -6, -18, 4, 5, -16, -20, -25, 23, 20, 33, 43, 40, 4, 34, 19, 20, 10, -17, 50, 54, -1, 17, 12, 10, -6, 7, -1, -2, -5, 3, -19, -6, -24, -41, -26, -44, -2, 45, 11, 2, 11, 21, 21, 31, 37, 37, 36, 53, -6, 13, -8, -8, -13, -18, -7, 16, 7, 18, -18, -16, -6, -64, -65, -29, 12, 12, -11, -14, 1, 54, 16, 6, -14, 53, 38, 56, 6, -11, 24, 15, -14, -19, 15, 8, 4, -1, 16, -5, 29, -15, -24, -3, -19, -21, -49, -59, 1, 18, 12, -5, -28, 15, -16, -7, -62, -59, -24, -14, 8, 1, -15, -21, 13, -13, 11, 6, -51, -30, -16, -9, -10, -53, -27, -44, -10, 64, 34, -25, -47, 2, 24, 2, -54, -72, -46, -31, 17, -4, -7, 14, -6, -16, -14, 11, -64, -31, -8, -5, -9, -52, -53, -43, 3, 62, 12, 6, -20, 1, -7, -4, -55, -52, -14, -49, -2, 20, 7, 6, 1, -9, -18, -40, -44, -41, 8, 3, -8, -29, -23, -29, 32, 53, -15, -2, 6, -16, -21, -30, -50, -36, -44, -30, -8, -17, -13, 17, 9, -4, -16, -36, -21, 12, -12, -15, -16, -41, 16, 21, 32, 59, -8, -10, 3, -50, -8, -17, -33, -59, -62, -23, -10, -8, -6, -18, -6, -2, -40, -7, -17, 17, -21, -79, -75, 4, 62, 47, 11, -3, -3, 11, -13, -34, 10, 4, -39, -42, -28, -23, -3, 8, -1, 6, 10, 17, -11, -51, -46, 0, -15, -31, -28, 3, 27, 17, -24, -14, -22, 10, -19, -13, 6, 17, -10, -40, -42, -37, -9, -7, -14, -16, 9, 15, -41, -59, -53, -16, -10, -3, -8, 4, 26, 24, -52, -29, -5, 3, -8, 22, 41, 17, 39, -49, -17, -15, 3, 16, -17, -20, -17, -18, 2, -14, -58, -24, -5, -24, 50, 63, 11, -19, -46, -26, 4, 15, 2, 1, 5, 12, 34, -27, -13, 2, -5, 8, 11, -11, 26, -32, -16, -11, -69, -29, -28, -59, 15, 50, -2, 8, -29, -47, 7, -10, 10, -25, -17, 6, 6, -31, -53, -27, -2, -15, 3, 10, -27, 25, 21, -30, -10, -11, -25, 20, 23, 4, 2, -13, -9, -33, -40, 10, 4, -8, 3, 8, 29, 9, -13, -16, 7, 14, -1, 4, -9, -6, -11, -17, -21, -15, -30, 41, 34, 23, 16, 12, -54, -6, -18, -65, -37, -27, -39, 22, 24, 3, -15, 16, 10, -5, -6, 1, -28, -15, 2, 14, -23, -34, 35, 70, 38, 29, 26, 11, -36, -36, -61, -32, -29, -45, -34, 32, 15, 35, -2, -23, 15, -15, 20, 14, 2, 18, 15, 16, 7, -15, 65, 82, 52, 13, -12, -3, -9, 12, -37, -53, -47, -29, -7, 28, 54, -4, 24, -2, 0, 9, -6, -12, -41, 13, 39, 49, -1, 20, 48, 70, 49, 5, 16, 10, 8, 22, -1, -56, -74, -75, -29, 49, 67, 47, 39, 22, 7, -15, 3, -14, -12, -7, 8, 57, 30, 32, 49, 50, 62, 8, 17, 11, 45, 2, -28, -58, -80, -52, -19, 23, 62, 68, 24, 22, 10, -3, -6, 18, -18, -14, -10, 41, 62, 42, 37, 43, 31, -16, -6, 33, 16, 5, -41, -53, -46, -74, -12, 5, 38, 48, 8, 5, 5, -2, -11, -20, 9, -20, -33, 13, 44, 59, 48, 59, 1, -17, -41, -19, -19, -17, 10, -49, -18, -44, -36, -57, 19, 62, 22, 8, -14, -19, 17, -4, 16, 15, -16, -25, 9, 30, 69, 44, 39, -26, -18, -43, -30, 9, 11, 7, -20, -25, -51, -10, -2, -9, -22, 13, -19, -5, 11, -10, -8, -19, -8, -40, 12, 20, 38, 3, 24, -20, -8, -21, 12, -4, 48, -4, -8, 2, -13, 9, 7, 21, 22, -9),
  86 => (4, 1, 14, -9, -18, -9, -1, -1, -18, -5, -10, 1, -5, 13, -9, -3, -23, -1, -10, 18, -18, -2, 9, -12, -4, -18, 12, 19, 1, -4, -5, -13, 19, -8, -2, 8, -4, -18, 15, -10, 20, -16, -14, -45, -44, -23, 31, 28, -6, 20, -13, -7, -16, -11, -7, 0, -9, -2, -1, -11, 12, -20, 13, 19, -17, -5, -41, -12, -20, 19, 27, -1, -67, -66, -39, 36, 19, 15, 31, -19, 7, -20, 18, -16, 8, -10, -2, -19, 4, 0, 8, 13, -19, 3, 13, -14, 11, -12, 0, -10, -8, 0, -26, -5, -11, -17, 21, 10, 5, -3, 15, -6, 11, -20, -6, -15, 16, -16, 14, 13, 12, -26, 16, 3, 0, -25, -23, 16, -8, -6, -32, -58, -34, 4, 13, 26, 10, -1, -3, 12, -3, 10, 17, 18, 0, -7, 0, 20, -13, 8, -11, -51, -33, 4, 44, 21, 17, -7, -64, -60, -2, -29, -14, 0, 16, -41, -20, -3, -12, -14, 14, 0, 0, -9, -14, -1, -6, 0, -11, -65, -59, -20, 20, 1, 21, 14, -41, -34, -7, -9, -30, 41, 14, -4, -2, 4, 7, -8, 2, -11, -19, 4, 26, -36, 41, 8, -26, -57, -55, -1, -6, 25, 15, 15, -10, -54, -21, 6, -3, 42, 25, 14, -21, -9, -2, -4, 4, -1, -11, -17, -11, -18, 16, -36, -24, -56, -24, -24, 5, 33, 19, 29, -25, -64, -16, -8, -26, -1, 53, 19, -52, -8, 7, -10, -7, 15, 1, 3, 14, -50, -20, 0, 12, -52, -54, -25, 28, 47, 9, 22, -12, -49, -35, -8, -29, 2, 44, 13, 5, -21, 5, 0, -5, 5, -8, 19, 30, 1, 17, 10, -4, -49, -44, -28, 24, 37, 27, 23, 14, -21, -30, -43, -26, 27, 18, 39, 8, -27, 21, -14, 6, 4, 3, 10, 54, 28, 17, -15, -5, -46, -60, -35, 3, 7, 4, 22, -44, -64, -59, -40, -64, -11, 17, 31, 42, 2, -12, -19, 20, 13, -4, 5, 62, 19, 20, 12, -1, -34, -45, -32, 7, 15, -3, 3, -33, -82, -29, -23, -7, 12, 28, 38, 10, -34, 4, -1, -9, 14, 20, 30, 74, 34, 19, 39, 14, -84, -81, -42, 21, 19, 21, 9, -20, -66, -82, -23, -8, -5, 13, 34, 12, -19, 9, 4, 18, 17, 3, 45, 59, 25, 38, 39, -32, -102, -65, -16, -21, 20, 14, 8, -10, -25, -96, -51, -15, -9, 20, 28, 32, 5, -13, 19, 5, -19, 22, 34, 62, 16, 15, 66, -26, -51, -70, -67, -25, 4, 0, 15, 15, -19, -69, -65, -19, 21, 39, 12, -1, 17, 15, -4, -11, 1, -1, 27, 48, 29, 44, 40, -26, -66, -43, -23, -18, 12, 21, -1, 5, -24, -67, -54, -26, -11, 47, 9, 23, 0, 7, -15, 9, -14, 10, 24, 14, 15, 29, 9, 8, -37, -54, -36, -8, 22, 28, 15, 45, -20, -49, -47, -47, -11, 26, 13, 32, 1, -16, 18, 6, 10, 11, 8, -5, -10, 36, 11, 16, -42, -66, -34, -20, 16, -8, 14, 19, 13, -71, -13, -45, -31, 1, 20, 62, 21, -16, 13, 14, -3, -36, 14, 1, 28, 3, 27, 43, -8, -58, -42, -4, 0, 19, 22, 16, -9, -37, -29, -47, -20, 10, 16, 17, 21, 0, 19, -1, 14, -42, 29, 26, 17, 29, 36, 50, -16, -32, -12, -29, -9, 17, 7, -10, 2, -52, -50, -45, -35, -5, 11, 27, -29, 8, -7, -4, 20, 13, 22, 54, 15, 15, 25, 27, -3, -17, -24, -34, 0, -19, 8, -12, -5, -9, -33, -50, -22, 12, 13, 3, -39, -16, -14, -15, -11, 21, 45, 39, 58, 30, 18, 21, 17, 8, -63, -20, 17, -8, 15, 20, -2, 4, 27, 7, -18, -1, 14, 11, -43, 18, 13, 12, 0, 8, -4, 22, 41, 8, 30, 30, 33, 5, -29, -14, 5, -22, 14, 18, 5, -1, -11, 1, -8, 17, 25, -21, -59, 14, 7, -8, -8, -12, 5, 15, 0, 26, -17, 7, 5, -10, -26, -27, 13, -5, -7, 11, 21, -12, -21, -10, 37, 28, -2, -5, 8, 8, -17, 8, 2, 39, 32, 6, 23, 13, 35, 16, -13, -11, -12, 2, -11, -28, -1, -14, 24, 9, 1, -28, 8, 45, 24, -6, -18, 13, 20, 10, -2, 6, 24, 1, -10, 20, 22, 48, 19, -2, 2, -16, -3, 3, 2, 1, 10, 26, -9, -2, 33, 34, 1, -16, 6, -17, -1, -14, 3, 10, 6, 0, -37, 23, 27, 28, 19, 18, -22, -26, -33, 12, 42, -6, -8, -23, 4, 20, 25, 7, 23, -11, -33),
  87 => (12, -1, 17, 4, 12, -3, 18, -16, 14, 6, -11, -13, 10, 0, 33, 19, -10, 26, 3, 26, 25, 15, 32, 15, -17, -5, -4, -17, -8, 19, 11, 9, -9, 10, 15, 1, -3, 15, -43, -26, -22, -6, -31, 11, 42, 47, 30, 50, 31, 64, 39, -3, 4, -20, -11, -12, -9, 0, 4, 16, 12, 0, -11, 7, 13, -39, -7, -10, -1, 67, 70, 62, 26, 33, -16, 35, 21, 18, 22, 16, -47, -12, -4, 9, -6, 9, -12, 15, 11, -14, 2, -2, 20, 7, -55, -23, 0, 22, 52, 43, 34, 35, 24, 26, 12, -17, -1, 16, -20, -25, -14, -20, 0, 0, -10, 14, -6, 11, -4, 34, -15, -62, -19, -34, -21, 25, 22, 10, 55, 21, 27, -2, -2, 49, 31, 35, -22, -33, -16, 8, -17, 10, 16, 14, 3, 12, 26, 40, 24, 24, 31, 11, -9, 9, 26, 11, 15, 0, 16, -23, -12, 32, 25, 41, -12, -25, 3, 8, 18, -2, -17, 15, 14, 4, 27, 57, -12, 32, 32, -5, -17, 27, 21, 8, 20, 47, -3, 10, -23, -23, 41, 38, 21, -2, 1, -5, -2, 4, 9, 21, 1, 12, 57, 34, 25, 59, 30, 0, 32, 66, 66, 62, 43, 36, 25, 29, 29, 19, 17, 29, -15, -13, 33, 40, -20, -7, 5, -2, 20, -5, 57, 66, 79, 56, 64, 47, 107, 119, 135, 109, 41, 13, 40, 29, -22, 0, -16, 17, 8, 29, 54, 59, -17, -3, -15, -18, 19, 12, 25, 42, 35, 49, 39, 55, 70, 111, 107, 68, 9, -33, 26, 29, 3, 32, 27, -12, -9, -1, 26, 21, 4, -17, 20, 14, -6, -6, 3, 12, 27, 34, 31, -9, 4, 45, 40, 25, 44, 24, 45, 36, 37, 8, 17, 11, 18, 15, -15, -7, -9, -18, 17, 15, 2, -68, -6, -34, 37, 28, 35, -2, -9, 0, 37, 47, 33, 2, 20, 16, 3, 12, 30, 31, -4, 1, 14, -4, -7, 11, 7, -15, 46, -47, 53, 35, 20, 18, 26, -6, -12, -19, 24, 26, 40, 40, 21, 9, 9, 19, 33, 54, 8, 46, 2, 33, -10, 10, -13, -12, 15, -52, 13, 58, 16, 18, 16, -10, -39, 24, 48, -2, 35, 55, 48, 11, -18, -4, 27, 46, 53, 71, 69, 64, -1, -4, 16, 14, 8, -20, 84, 59, 52, 37, 65, 35, 29, 12, 19, 35, 30, 30, 34, -8, 4, 18, 20, 49, 50, 81, 46, -20, 16, 16, -10, -12, 38, 50, 115, 41, 34, 4, 16, 27, 12, 55, 47, 37, 43, 39, 27, 9, 30, 13, 55, 54, 40, 53, 15, -4, -11, -7, 7, -3, 19, 17, 50, 7, 35, 10, -26, -6, -18, 32, 14, -5, 37, 38, 58, 16, -14, 39, 42, 58, 16, 31, 21, -26, 0, 15, -12, -12, -1, 46, 12, -12, -11, -3, -8, -28, 29, 5, 20, 19, -6, -4, 42, 1, -11, 13, 21, 53, 15, 8, -33, -38, -15, 12, -12, -12, 6, 25, -6, -21, 12, -35, -32, -3, 10, -2, -16, 14, -2, 1, 13, -1, 4, 26, 1, 0, -7, 5, -20, -55, -19, 0, 14, -4, -6, 35, 9, -10, -14, -22, 14, 21, -24, -15, -4, -9, -1, 17, 33, 10, 7, 18, 9, -5, -19, 19, 1, 5, -6, -21, 19, 20, -17, -1, 15, -8, 7, -11, 3, -14, -24, 12, 27, -38, -19, 1, -18, 23, -37, -74, -37, -4, -12, -19, 3, -10, -7, 15, -3, 4, -18, 6, 15, 12, -2, 25, -1, 0, 11, -13, 26, -14, -34, 31, -24, -26, -53, -62, -9, 4, -41, -41, -28, -45, -3, -8, -18, 17, -34, 14, 34, 14, 20, 14, -10, -19, -16, -32, -30, 3, -25, -1, -22, -8, -28, -49, -13, 10, 33, 18, -36, -78, -14, -1, 20, -3, -10, 22, 20, 22, 25, 18, -51, -26, -14, -34, -34, -14, -20, 0, 8, -1, 5, 2, 16, -4, 64, 11, 11, -30, -11, 11, 5, -3, -43, 53, 16, 55, 62, 16, -5, -22, -4, -20, 14, -8, -22, 0, 25, 18, -6, 6, -12, 20, 35, 43, 9, 4, 13, 10, 16, -5, 2, 1, 47, 55, 39, 60, 15, 14, 23, 15, 35, 29, 12, 45, 20, 21, -26, -10, 13, 20, 35, 62, 3, 0, 5, 8, -19, 7, 24, 38, 50, 46, 34, 57, 42, 61, 53, 40, 45, 22, 72, 50, 45, 29, 18, 23, 29, 60, 26, 20, -18, 2, 0, 11, 19, -10, -7, 35, 33, 49, 35, 29, 63, 76, 78, 44, 69, 31, 84, 104, 98, 49, 18, 14, 58, 37, 16, 13, -50, -32),
  88 => (6, 17, -2, 4, 19, -18, -16, 4, 13, 6, 18, -20, -6, -8, 35, 35, 10, -23, -47, -19, -18, -4, -19, 0, -16, -16, -18, -8, -14, 19, 14, -17, -14, 16, 10, -13, -4, -10, -28, -25, 32, 52, -3, 41, 2, -8, -22, -1, 24, 50, 2, -15, -2, -9, -2, -13, -6, -4, 6, 20, -1, 1, -3, 6, -18, -22, 13, 21, 45, 24, 3, -40, -35, -46, -21, -10, -12, 6, 48, 5, -38, -45, 13, 6, 3, 8, 1, -17, 15, 16, 5, 1, -11, 6, -4, 12, -12, -20, -45, -25, -14, -14, -5, 17, -14, 18, 13, 15, 34, -22, -6, 20, 20, -15, -1, -19, 10, -19, -7, 1, -19, 36, 31, 7, 0, -17, -20, -26, -27, -17, -37, 20, 25, 2, 6, -4, 48, -37, -11, -11, 0, 20, -15, -16, 7, 5, -3, 7, 32, 68, 35, 8, 2, 7, 29, 33, 1, 14, 38, 39, 41, 37, -6, 36, 40, -5, 15, 5, 11, 0, 12, 12, 6, 16, 1, 16, 87, 96, 69, 49, 73, 44, 26, -10, 0, 22, 21, 51, 51, 66, 24, 9, 9, 8, -30, 2, -7, 1, 11, -20, -10, -3, 9, 47, 108, 116, 94, 75, 64, 20, 17, 4, -18, -10, 7, 12, 44, 19, 67, 21, -39, 9, -20, 42, 14, 16, 0, -14, 2, 5, 43, 89, 103, 114, 102, 73, 47, 25, 49, 42, 44, 45, 40, 98, 26, 34, 27, 60, 1, 5, -8, 72, 5, -7, 9, -14, -11, 6, 64, 95, 81, 33, 5, 50, 37, 26, 70, 39, 13, 44, 26, 59, 29, 0, 32, 42, -19, 23, 21, 60, -3, 18, 7, -13, -7, 37, 93, 60, 40, -11, -22, 41, 38, 31, 24, 46, 13, 26, -12, 30, -4, -51, -27, -15, -2, 14, 2, 36, 19, 15, 17, -3, -1, 61, 38, 26, 46, -10, 10, 40, 45, 44, 23, 26, 5, 30, -10, -27, -15, -18, 19, -10, -9, -30, -31, 18, -5, 3, -16, 0, -7, 17, 14, 10, 8, -38, 15, 45, 47, 20, -6, 3, 12, 5, 19, 18, -2, -4, 9, 11, -19, -54, -60, 8, -12, 2, -5, -17, -4, 21, -41, -23, -16, -6, 42, 61, 29, -7, -6, 18, 49, 26, 25, -1, -3, -14, -42, -35, -61, -97, -54, -1, 10, 14, 6, -19, 14, 8, -16, -28, -4, -6, -8, 5, -12, -48, -39, -14, -6, -9, 8, 5, -23, -9, -31, -40, -40, -62, -55, 7, -1, 3, 5, -7, 12, -11, 9, -53, -70, -74, -106, -97, -66, -55, -34, 8, 0, 9, 13, 10, -21, -38, -9, -38, 13, -34, -22, 61, -10, -10, -8, 9, -46, -16, -68, -57, -73, -96, -107, -65, -54, -25, -30, 6, 12, 28, 45, -23, -26, -2, -19, -23, -7, -5, 6, 37, 4, -1, 11, -12, -57, -33, -67, -38, -64, -64, -44, -46, -7, -32, -8, 6, 36, 21, 0, -6, -17, 14, -27, -30, -40, -66, -9, 54, 6, -7, -6, 11, -79, -17, -18, 5, -37, -27, -34, -20, -9, -26, -9, -1, 26, 11, 17, -15, -28, -11, -9, -47, -6, -52, 20, 70, -3, -9, 21, 20, -14, 9, 12, -5, 0, -6, -26, -5, -12, -58, 16, 29, 35, 6, 8, -28, -33, -27, -30, -28, -32, -29, 17, 69, 1, 12, -11, 7, -39, 7, 9, -10, -32, -8, -4, -14, -9, -15, 18, 34, 47, 16, -8, -43, -43, -12, -8, -64, -29, -13, 10, 51, 13, 10, 4, -17, 18, 19, 1, -9, -3, 24, 50, 25, -6, 16, 13, 32, 35, 29, -1, -5, -5, 28, -29, -43, -24, -24, -23, 3, 8, 3, 8, -9, -9, 55, 21, -31, -29, 17, 38, 1, -8, -9, -15, 28, 50, 16, 11, -14, 25, 54, 18, 2, -53, -21, -38, -22, 15, 2, 15, -12, 11, 29, 27, -34, -61, 3, -1, -4, -5, -22, -1, 11, 10, 22, 16, 19, -6, 31, -2, -13, -44, -26, -80, 3, 17, -17, -11, -17, -11, 25, 11, -7, -34, 25, 0, -23, 12, 3, -9, 9, 5, 17, 17, 39, -14, 35, 18, -18, -28, 5, -7, 1, -2, -17, -7, -7, 29, 49, 47, 4, -27, 17, 28, 7, -1, 19, 16, 30, 39, 14, 6, 2, -1, -14, -3, 4, -20, 11, 15, 14, 1, -9, 10, -16, 24, 57, 62, 25, -35, 8, 35, 11, -1, 28, 28, 40, 43, 30, 12, 3, -1, -11, 4, -12, 20, 18, 32, 22, -15, -10, -8, -5, -12, 4, 63, 47, 33, 3, 50, 43, 31, 42, 44, 65, 63, 72, 25, 27, 50, 53, 59, 85, 21, 50, 56, 4),
  89 => (-5, -10, 2, 8, 20, -2, 16, 6, -19, -12, 20, -12, 12, 8, 32, 0, -34, -24, 7, 31, 26, 5, -29, 3, -13, 8, 10, 7, -10, -10, -14, -2, -13, -20, 13, 12, 13, -10, 20, 46, 12, -9, 24, 10, 49, 48, 40, 54, 42, 79, 44, -13, -26, -5, 20, 1, -15, 9, 15, -7, -21, -17, -7, -4, -19, 32, -12, 40, 29, 3, 18, 51, 46, 45, 55, 21, -9, -22, -32, -34, -46, -11, 7, -4, 19, 9, -12, -3, -5, -13, 8, 3, 6, 3, 40, 0, -7, 41, 54, 37, 40, 7, 19, 43, 6, -16, 14, -2, -1, -13, 11, -17, -5, -3, -13, -9, -11, -17, 6, -7, -1, -20, -6, -15, -28, -3, -3, 38, 25, 7, 28, 22, -2, -3, -1, 13, 43, 10, -10, -10, -1, 16, 20, 15, -14, -8, 8, 29, -54, -43, -48, -68, 3, 8, 19, 31, 32, 53, 26, -8, -8, 13, 21, 39, 50, -28, -16, 15, -18, 1, 8, 18, 11, -13, 25, 33, -35, 30, -21, 8, 38, 31, 33, 47, 39, 15, 16, 43, 38, 28, 49, 45, 34, -31, 1, -2, 3, 2, -9, -17, 10, 0, 50, 47, 42, 49, 48, 44, 9, 27, -2, 42, 21, 2, 10, 7, 4, 30, 38, 31, 34, -9, 35, -7, 20, 3, -9, 7, 3, 5, 54, 46, 42, 32, 44, 11, -5, 20, 13, 21, 17, 20, 4, 4, 28, 38, 45, 14, -11, 3, 32, 25, 2, 2, -8, -17, 0, -15, 43, 47, 36, 51, 28, -11, -13, 0, 33, 56, 53, 10, 41, 40, 17, 10, 18, 8, -14, 8, -20, -1, 12, 6, 0, -4, -3, -26, 74, 70, 68, 78, 42, 9, 19, 29, 49, 66, 20, 5, 32, 12, -15, -15, -24, -30, -30, -14, -6, -7, 8, 12, -16, 16, 0, -21, 45, 51, 42, 70, 27, 15, -3, 41, 2, 47, 40, 19, 24, 1, -17, -41, -32, 10, 6, -21, -20, -26, 10, -17, 11, 3, 3, -19, 50, 22, 29, 26, 2, 4, -45, 15, -23, 25, 39, 10, 21, -25, -24, -12, -5, -2, 20, -31, -28, -62, -11, 1, -10, 13, 8, -25, 29, -34, -15, -53, -38, -87, -32, -54, -33, -2, 7, -11, -17, 3, -10, -7, -10, 6, 1, -50, -21, -3, -12, 0, 10, 20, 17, -7, 4, -41, -54, -66, -46, -70, -69, -74, -69, -73, -47, -8, -2, -8, -31, -56, 4, 7, 20, -25, -13, -30, 11, 15, 4, 19, 22, -14, -14, -42, -51, -45, -16, -43, -59, -29, -47, -36, -31, -10, -50, -22, -41, -42, 29, 22, 8, 32, -32, -64, -8, 18, -11, 6, -9, -20, -18, -30, 3, 28, 1, -10, -5, 5, 31, -19, -31, -50, -61, -32, -16, -13, 36, 27, -6, 65, -6, -30, 3, 19, -9, 1, -30, -5, -7, -5, 39, 10, 21, 62, 25, -16, -5, -14, -42, -28, -22, 5, 10, 8, 5, 12, 28, 51, 44, -44, 0, 15, 5, 5, 2, -28, -15, -29, -22, 21, 40, 47, 19, -11, -33, -8, -28, -25, 1, -16, -8, -9, -1, 17, -2, 28, 69, 8, 4, -17, -5, -14, -15, -42, 5, -17, -30, 16, 39, 64, 19, 15, 32, 6, -18, 17, 28, 18, 46, 42, 11, 39, 21, 34, 29, -35, -10, 5, 19, 12, -3, -32, 7, 17, -10, 19, 63, 45, 55, 41, 30, 43, 28, 58, 50, 33, 40, 8, 16, 37, -2, 20, 46, -9, -3, 19, -14, 2, -27, 10, 6, 1, 14, 22, 44, 53, 44, 50, 32, 47, 50, 48, 65, 63, 60, 27, 16, 19, 19, 10, 63, 25, 11, -18, 0, -8, 4, 19, 11, 34, 26, 39, 45, 47, 43, 39, 46, 23, 50, 39, 68, 85, 69, 19, -25, 23, 1, 25, 70, 26, -13, 3, 21, -4, 10, 23, 55, 49, 61, 47, 69, 48, 39, 31, 16, 33, 60, 33, 56, 57, 44, -3, 5, 39, 29, 17, 39, 6, -8, -3, -4, -5, 3, 27, 35, 40, 18, 37, 60, 22, 8, -2, 23, 18, 71, 52, 67, 53, 33, 18, 36, 68, 19, 13, 5, 1, -19, 13, 17, -10, -26, 9, 52, 24, 22, 35, 33, 30, 36, 27, -3, 27, 56, 27, 30, 41, 22, -11, 0, -6, 10, -11, -6, 44, -13, 17, -20, -13, -13, 46, 34, 26, 43, 46, 51, 58, 37, 11, -15, -28, -49, -39, -20, 8, 14, -16, 30, -17, -17, -4, 24, 9, 16, 17, -6, -10, 10, 9, 42, 53, 14, 42, 46, -10, -17, -7, -33, -34, -18, -39, -13, -8, 34, 11, 52, 12, 47, 1, -17, 8),
  90 => (-3, -13, 6, -15, -5, -13, -10, -13, -15, 20, -4, 18, -12, -20, 15, 17, 1, -19, -9, 7, -40, 5, 13, 11, -13, 8, -13, 19, -20, 9, 4, -17, -1, 18, 20, -17, -20, 15, -16, 8, 21, 4, 18, -13, 14, 0, 5, 8, -18, -28, 17, -19, -15, 8, -6, -3, -14, 15, -4, 4, 14, -12, -4, 12, -13, 1, 45, 38, 25, 22, 6, 27, 16, 15, -22, 1, 19, 30, 35, 46, -1, -22, 16, -5, 17, 1, 16, 15, 19, -11, -9, -19, -6, -3, 4, 5, -8, -19, 10, -8, 5, -18, -27, 11, 10, 54, 56, 41, 30, 14, -9, -10, -14, 1, -13, -10, 15, -20, -12, 10, -1, 18, 4, 2, -13, 10, -23, -24, -18, 3, -2, 17, 24, 37, 25, 6, 14, 15, 7, -19, -5, 16, 6, -12, -3, -2, 26, -2, 10, 3, 0, 8, -12, 13, 2, -7, -1, 11, -2, 23, 33, 16, -4, -31, -38, 16, -1, 6, -8, 13, 12, -6, -6, 20, 30, -9, -2, 1, 3, -17, -38, 19, -27, -41, -35, -21, -44, -10, -19, -42, -52, -49, -22, -24, 11, -4, 1, -4, -5, 8, -1, 19, 31, 3, -10, 19, 14, -19, -22, -40, -90, -98, -89, -129, -113, -67, -101, -124, -134, -132, -29, -7, -34, -8, 12, 9, -3, -3, -17, 4, -7, 54, 14, 33, 35, 33, 21, 35, 3, -3, -21, -29, -3, -14, -19, -16, -65, -52, 3, -45, -10, -31, 13, -2, 6, 7, -20, -15, -11, 48, 19, 65, 28, 52, 37, 53, 25, 5, 13, 19, 15, 44, 23, 27, 26, 44, 25, -1, -32, -46, 9, -1, 2, 0, -9, -10, 0, 22, 17, 19, 7, 4, 18, 37, 39, -4, 3, 6, 5, 28, 42, 74, 55, 58, 76, 19, -15, -30, -9, 10, 19, -7, -11, -3, -2, -9, -19, -32, -62, -45, -40, -11, 33, 26, 36, 40, 76, 73, 98, 66, 43, 29, 33, 18, 33, -12, -12, 19, -19, 7, 11, -4, -24, -17, -31, -77, -4, -24, -69, -43, -70, -41, -4, 7, -9, 2, 7, -6, -10, -9, 15, 39, 43, -4, -19, 9, -12, -6, -3, -28, 3, 0, -1, 5, 7, -30, -20, -65, -50, -53, -40, -65, -63, -81, -81, -92, -71, -49, -26, -2, 69, -14, -3, 11, 12, -1, 27, -2, -15, 13, 45, 36, 13, 9, 22, -14, 11, 3, -20, -53, -57, -81, -98, -82, -95, -81, -43, -16, 40, 7, 6, -6, -8, -7, -12, 13, 5, 10, 31, 49, 37, 2, 17, 16, 16, 22, 31, -1, 25, 8, -30, -22, -8, -46, -68, -27, 21, -18, 13, 1, 4, 17, -4, 5, -12, -8, 9, 7, 15, 20, 10, 5, -1, 6, 3, 9, 18, 32, 1, 30, 40, -26, -21, 6, 28, 2, -14, -18, -17, 5, 7, -15, -25, -17, 12, 10, 9, 0, 35, 17, 42, 6, 3, 0, 24, 6, -4, -14, 7, 20, -24, -57, -43, 14, -3, 3, 5, 12, -26, -48, -23, 2, 4, -47, -43, 8, 8, 14, 31, 23, -22, 9, 42, 4, 23, 13, -1, 15, 38, -64, -56, -8, 10, -5, 4, -4, -12, -39, 4, -3, -2, -39, -48, -16, -2, -38, -1, 21, -4, 14, 5, 20, 10, -6, -16, -10, 30, -18, -12, -30, -20, 2, 7, 6, -11, -30, -22, -42, -29, -27, -27, -25, -9, -19, 7, -1, -22, -23, -1, 7, 6, 4, -20, -14, -28, -55, -27, 20, 21, -16, -5, 2, 7, -48, -51, -36, -34, -37, -25, 8, -7, -21, -16, 18, -31, 9, 14, 3, -9, -6, 13, -59, -49, -51, -31, -33, 21, -20, -16, 13, -16, -16, -5, -55, -20, -18, -16, -4, -28, -9, 5, 9, -35, -14, -8, -37, -20, 17, 26, -25, -60, -29, -11, -72, -21, -8, -11, -9, 12, -24, -13, -17, -2, -31, -1, -5, 8, -6, 6, -8, -31, -6, -12, -31, -1, -8, 10, -28, 21, 8, -2, -39, 16, 6, 6, 12, -15, -45, -45, -21, 3, -17, -6, 12, -16, -6, -13, -34, -30, -22, -24, -21, -32, 1, -1, -9, 21, 29, 9, -10, -13, 13, 1, -8, -20, -29, -56, -50, 15, 19, 1, 11, 9, 17, -10, -29, -29, -3, -16, -5, 21, 10, 25, 9, -9, 14, 3, -14, 0, 18, 18, 0, -25, -12, -10, -15, -28, -27, 13, 28, 37, 4, -31, -6, -34, -14, -22, 4, 6, 30, 41, -2, 22, 25, 17, -11, -16, -6, 17, -17, 16, -2, -17, 7, 33, -17, -10, 14, 38, 29, 23, -8, 14, 7, 25, 34, 33, 59, 46, 28, 52, 15, 10, -14),
  91 => (-9, 2, -20, 2, 9, -12, 5, 6, -11, -20, 14, -14, 13, -19, -30, -26, -56, -8, 0, 29, -6, -13, 7, -4, 13, 19, 20, 20, 4, -2, 20, -12, 18, -5, 3, -8, 8, 11, -17, 13, -8, -11, -35, -16, -25, 4, -20, -31, -32, -18, -27, -16, -15, -14, 10, 9, 8, 21, 8, -10, -14, -2, 9, -4, 11, 5, 12, 5, -5, -14, -25, 19, 21, 15, -2, -16, -21, 21, 22, 7, 3, -8, -4, -1, -15, -12, -5, -1, 8, 2, -8, 10, -7, -9, -25, -20, -71, -12, 1, 39, 62, -10, 6, 2, 21, -4, 0, 11, -41, 28, -5, -3, 5, 0, -2, -17, -5, -14, -12, -36, -21, -34, -78, -75, -37, -8, 48, 46, 16, -16, 5, 6, 18, -24, -41, -59, -32, -14, 5, -3, 17, 12, 1, 14, 3, -14, -53, 29, -28, -103, -141, -75, -3, 17, 35, 42, 31, 9, 16, -1, -23, -46, -21, -67, -84, -25, -15, 9, -13, -12, 18, -1, 16, -18, -53, 56, -26, -83, -114, -15, 37, 25, 18, 12, 23, -6, -10, -37, -68, -85, -36, -23, -42, 6, 13, 13, -14, -4, 9, -10, -2, 8, 11, -9, -3, -100, -57, 29, 41, -7, 33, -3, 12, -52, -59, -26, -34, -86, -58, -31, -17, 12, -16, -21, -18, -11, 10, 14, -20, 11, 19, -4, 8, -49, -34, 34, 12, 33, 16, 1, -13, -80, -103, -34, -11, -58, -78, -39, -9, 28, 1, 18, -8, -7, -10, 3, 11, -21, 12, 51, 8, -41, 26, 10, 40, 13, 5, -10, -16, -74, -50, -24, -16, -45, -5, -3, 12, 35, -12, 19, 2, -9, 1, 20, -20, 18, -16, 13, -34, -26, -45, 9, 23, -12, -23, -46, -20, -29, -34, -11, -5, 4, -13, 49, 18, 18, 3, -19, 18, -17, 14, 20, 0, 19, -5, 4, -20, -38, -8, 26, -27, -41, -41, -5, -10, -37, -21, -3, 27, 23, 14, 27, 53, 8, 27, -38, 3, -15, 17, 9, 18, 16, 24, 13, -24, 11, 41, -12, -8, -7, 3, -18, -28, -14, 18, 8, 12, 38, 54, 38, 28, 25, 15, -12, 8, 8, -14, -12, 29, -12, -36, 10, 24, 18, 36, 7, -17, 17, 12, 28, 11, 14, 18, 16, 20, 43, 34, 52, 59, 35, 36, -46, -13, -9, 18, 2, 1, -61, -31, -2, -17, -11, 25, 3, 4, 33, 35, 20, 52, 15, 4, 38, 31, 16, 26, 22, 31, 2, 23, -9, 11, 7, -13, 16, -20, -32, -18, 21, -14, -14, 21, 6, 25, 26, 54, 31, 44, 34, 10, -2, 20, 6, 27, 25, 2, -14, 3, 37, 20, -20, 7, 3, -18, -16, -18, 29, -6, 9, 14, -1, 26, 16, 11, 20, 10, 15, -9, 4, 9, 12, 23, 11, -7, -38, 6, 23, 19, 6, -11, 1, -13, -7, -8, -9, 1, 30, 14, -32, 43, 42, 16, 4, -7, -24, 8, 31, 32, 24, 16, 1, -22, -40, -15, 23, 3, 5, 3, 14, 25, 42, 30, -1, 0, 35, 14, -9, 0, 27, 36, 24, 14, 15, -1, 20, 7, -26, -10, -24, -40, -54, -75, -36, -10, -2, 12, -6, 51, 4, -5, 2, 31, 43, -16, -31, -14, -26, -7, 3, -11, -12, -23, -12, -31, -14, -15, -21, -31, -77, -81, -31, -10, 1, 14, -10, 10, -21, 1, -18, 0, 24, -32, -16, -20, -77, -64, -63, -96, -98, -66, -71, -36, -88, -45, -36, -69, -73, -54, -64, -1, -10, 19, 3, 20, -10, -10, -31, -15, 39, -6, -62, -70, -72, -68, -80, -91, -98, -71, -71, -85, -93, -45, -18, -96, -45, -60, -42, -14, 17, 11, -13, 19, -15, -17, -13, -3, 31, 2, 20, -33, -45, -57, -65, -89, -66, -66, -37, -62, -80, -77, -74, -45, -51, -45, -62, 8, -11, -3, 15, 9, 27, -4, 16, 10, 12, 5, 46, 7, -8, -68, -75, -85, -74, -32, -30, -8, -50, -38, -36, -42, -52, -18, -5, -2, -9, -4, -19, 8, -2, 31, 8, -19, -8, -21, 41, -29, -10, -21, -61, -96, -44, -42, 9, -5, -18, -42, -55, -75, -30, 9, -6, -20, 16, 0, 1, 3, 20, 12, 13, -34, -30, -49, 17, -35, -28, -25, 0, -16, -46, -37, 10, -15, -36, -22, -48, -34, -32, -21, -14, 1, 3, -8, 2, -18, -18, 4, -18, 8, -27, -50, -28, -6, -26, -17, 14, -27, -24, -21, -35, -33, -19, -6, -19, -13, -15, -16, -24, -8, -15, -15, -5, -8, -20, 0, 5, 5, 20, -16, -20, -33, -33, -4, -8, -5, -25, -16, -27, -18, -16, -23, -28, 20, 11, -3, -11),
  92 => (-16, -19, -2, -13, -1, -16, 1, -6, -13, 9, -7, 20, 11, 2, 18, 1, -14, 1, -1, 11, -14, 0, 4, -17, 15, 16, -3, 6, 12, 12, -20, 8, -15, 21, 3, 3, 12, -5, -18, -14, -9, -38, -57, -86, -70, -58, -22, -7, -39, -22, 8, 4, -21, 9, 0, 13, 13, -14, 4, 9, 11, -8, -5, -10, 8, 9, -11, -27, -35, -37, -22, 26, 10, 34, 36, 32, 18, -1, -28, -15, -11, -5, 13, -20, -1, -10, 1, -6, -20, -18, 13, 9, -7, 22, 30, 43, 36, 6, 6, 15, -2, 13, 28, 20, 20, -9, -31, -28, -13, 14, 4, 20, -7, -13, 3, 19, -10, 7, -12, 3, -42, 3, 50, 8, -1, -16, 12, 44, -4, 1, -27, 19, 38, 23, -9, -27, 3, -2, 12, 16, 7, -10, 5, -5, -12, 16, 22, 22, -33, 26, 6, -47, -20, 10, 18, -4, -29, -20, 19, 18, 21, 19, -7, -14, 25, -12, 11, 7, -1, -14, 17, 9, 10, 10, 29, -22, 28, 2, -69, -85, -9, 45, 21, 17, 29, 37, 7, 26, 4, 12, 2, 4, 10, -2, 0, -2, 4, 18, 15, 9, -21, -1, -21, -7, -9, -15, -43, -25, 13, 46, 12, 39, -2, 11, 47, 42, 16, -3, -22, 1, 19, 39, -7, -5, 18, -7, -16, 18, 6, 4, 10, 12, -67, -37, -14, 10, 28, 19, 30, 25, 15, 15, -3, 12, -18, -56, -78, -46, -26, 14, 3, 13, 11, 19, -19, -10, 10, 2, 41, -3, -90, -58, -36, -11, -3, 9, 30, 20, 18, 12, 2, -35, -70, -101, -87, -44, -23, -7, 1, -13, 6, 15, 8, 15, 15, -3, 23, 15, -52, -55, -39, -15, -10, 12, 3, -7, -6, 8, -37, -73, -74, -90, -59, -1, -29, 13, 13, -8, -10, 12, -8, 6, 1, -16, 24, -8, -41, -67, -26, 34, 17, 25, 11, -26, -15, -34, -49, -68, -70, -40, -51, -51, -16, -24, 14, 11, 2, 1, 15, 18, -8, -54, -3, -29, -51, -3, 29, 53, 60, 15, 14, -21, -1, -7, -46, -56, -74, -60, -63, -64, -59, -8, -7, -26, 4, -11, 4, -17, -12, -38, 2, -14, 8, 43, 48, 11, 7, -38, -63, -34, -23, 4, 10, -25, -40, -77, -83, -44, -23, -33, -2, -11, 19, -12, 19, 10, -21, 16, 7, 29, 31, 19, -5, -15, -49, -88, -19, -38, -45, 17, 22, 2, -79, -100, -78, -66, -35, -1, 1, -6, -12, -6, -1, 15, -48, -29, 9, 5, -14, 29, 31, -21, -31, -30, -42, -23, -1, 24, 22, -21, -79, -101, -52, -40, -14, -25, -11, -1, -4, 8, 11, -16, -72, -47, -30, -17, -21, 42, 59, 19, 1, -32, -40, -45, -33, 9, 20, -18, -82, -80, -65, 0, -8, -29, -4, -25, 18, -4, -16, -5, -67, -46, -40, -15, 6, 29, 43, 27, -15, -32, -34, -44, -44, -6, 25, -8, -45, -61, -11, 10, 0, -26, -2, 9, -17, -5, -4, 20, -68, -36, -47, 14, 39, 40, 26, 18, -1, -29, -48, -61, -31, -6, -11, 22, -26, -37, -12, 1, -35, -24, -33, 11, -12, -2, 15, 1, -34, -33, -43, 28, 76, 54, 33, 23, -2, -51, -65, -30, -25, 15, -1, 22, -22, -12, -18, -22, -51, -29, -13, 7, 1, 8, 11, -3, -19, -17, -24, 25, 59, 94, 52, 11, -2, -34, -33, -64, -60, -38, 10, 48, -6, -3, -31, -47, -48, -34, 7, -21, 1, 19, 5, -15, -43, -67, -22, 26, 72, 82, 19, 12, 5, -9, -20, -20, -41, -35, 25, 50, -5, -21, -47, -38, -18, -22, 10, -11, -5, -12, -20, 10, -23, -51, 42, 9, 1, 18, 12, -18, -20, -22, 8, 11, -8, -5, 9, 20, 18, -42, -23, -36, -3, 12, 14, -12, 11, -16, -10, 4, -5, -23, 2, -16, -26, -9, 4, -17, -15, -14, -27, -7, 11, 8, 7, 17, -26, -52, -67, -12, -27, 9, -2, 17, 11, -9, -7, 9, -43, -28, -28, -32, -23, 8, -5, -3, -1, -33, -22, -4, -1, -17, 18, -13, -28, -36, -15, -44, 20, 33, 14, -3, 10, 14, 18, -14, -34, -16, -31, -42, -28, 9, 30, 30, 31, 19, -4, 19, -2, 14, -12, -23, -62, -29, 3, -11, 9, 10, 1, -11, -3, -12, 5, 4, -27, -35, -11, -65, -40, -25, -28, -64, -43, -29, 8, 30, 22, 5, -24, -3, -36, -9, 5, -1, 6, 23, -11, 10, -14, 19, -6, -9, -8, -10, -33, -47, -29, -14, -37, -60, -16, 8, 18, 5, -15, -46, -75, -31, -2, 19, -22, -54, 12, 4, -4, 19),
  93 => (-4, 1, 15, -6, 7, -20, 18, -2, 5, -17, 0, 12, -18, -13, 22, 23, 14, 1, -50, -65, -43, -19, 1, -9, -19, -3, -15, -5, -20, 3, 6, 12, 16, -19, -20, 16, 4, 16, 31, 21, 35, 28, 17, 39, 30, 10, 14, 20, 27, 6, 47, -30, -25, -17, 4, 13, 1, -13, -15, -10, -20, 19, -9, 9, 20, 30, 45, 91, 37, 44, 38, 34, 21, 62, 37, 57, 61, 28, 10, 5, -71, 6, 5, -4, 10, 16, 12, -20, 2, 20, 13, -4, 17, 40, 36, 22, 25, 51, 34, 10, 44, 43, 53, 17, 28, 12, 49, 25, -63, -51, -8, 7, 14, 0, 7, 12, -6, -12, -7, 21, 56, 3, 1, -10, -23, -8, -2, 9, 64, 32, 50, 32, 33, 15, 45, 24, -25, -19, -20, -15, -18, -20, -17, -5, 6, 20, 47, 57, 17, -17, -3, -31, 8, 17, 31, 13, 12, 57, 42, 31, 12, 53, 5, 13, 54, 20, -18, -8, 5, 10, -9, -8, 4, 17, 10, 73, -15, 5, 26, 4, 15, 7, 14, -7, -9, 23, 10, 5, 45, 35, 13, 16, 59, 14, 24, 19, -13, 10, 1, 16, 17, 4, 47, 25, 42, 25, 15, 34, -4, 18, -4, 11, 2, 11, -8, 33, 48, 79, 66, 6, 36, 25, 38, 28, 19, -16, -18, 15, 20, 17, 16, 73, 53, 60, 65, 31, 26, 38, 26, 24, 8, 18, 35, 31, 26, 40, 42, 7, 52, 35, 24, 17, -11, -20, -18, 17, -16, -15, 64, 76, 58, 81, 54, 68, 76, 102, 109, 85, 30, 57, 57, 21, 35, 28, 50, 31, 44, 70, 8, 5, -11, -7, -1, -6, -20, -3, 49, 64, 66, 61, 52, 53, 70, 86, 90, 47, 22, 14, 21, 27, 17, 9, 3, 13, 16, 65, 61, 18, -12, -11, -15, -13, 2, -12, 48, 34, 79, 84, 64, 96, 70, 72, 61, 53, -26, -9, 7, -6, -12, -3, 12, 24, 33, 30, 50, 46, -11, -6, 12, 21, 29, -71, 35, -10, 46, 66, 53, 47, 77, 37, 27, 14, -11, -47, -33, -21, -23, -45, -5, 9, 22, 36, 7, 16, 11, -12, -6, -18, -13, -56, -9, -24, 32, 36, 20, 32, 39, 32, 38, 33, 7, -34, -25, -21, -7, -8, 3, 0, -4, -7, 9, 23, -15, -16, 7, 12, -28, -46, -29, -16, 6, -1, -22, -36, -5, 26, 20, 16, 26, -10, 11, -5, 7, -15, -4, -4, -2, 38, 17, 22, 9, -21, 18, -6, 7, -16, 20, 5, 11, -21, -35, 12, 7, 29, 34, 45, 42, 31, 19, 20, 5, -5, 10, 44, 41, 46, -6, 14, 17, 16, -3, -16, 36, 33, 15, 3, 33, 34, 3, -8, 38, 13, 36, 59, 48, -9, 25, 15, 20, 59, 4, 15, 30, 21, 36, 36, 5, -9, -17, 7, 7, 10, 48, 6, 5, -6, 5, 27, -4, 19, 5, 6, 24, 20, 0, 20, 44, 30, 27, 11, 68, 25, 61, 46, 9, -20, 9, -13, 33, 41, 29, -20, -25, -24, 21, -11, 19, 5, -17, 27, 22, 5, 12, 30, 48, 37, 24, 30, 39, 34, 89, 37, -9, 7, 6, 8, 10, 19, 52, 15, 11, 22, 36, 31, 13, 1, -4, 28, 19, 40, 21, 26, 41, 19, 10, 58, 12, 10, 32, 9, 16, -6, 19, 16, 2, -2, 12, 11, 18, 13, 23, -3, -20, -8, -13, -25, 38, 28, -15, 3, 54, 37, 58, 51, 60, 46, 40, 20, 9, -5, -1, 14, 28, -6, 7, 8, -4, -9, 32, 17, 28, -18, -7, 2, 15, 36, 12, 71, 65, 20, 56, 76, 73, 69, 45, 7, -20, 20, 16, -7, 29, -6, 28, 19, 2, -22, 9, 11, 39, 23, 28, 26, 26, 1, 22, 44, 54, 51, 31, 39, 56, 72, 22, 35, -8, -9, -1, -18, -9, 10, 49, 14, 8, -2, -16, -2, 0, -8, 9, 12, 46, -5, 24, 16, 39, 16, 45, 20, 17, 53, 41, 3, 6, 10, -18, 17, -17, -17, 12, 12, 25, 27, 22, 12, 26, 16, -5, -13, 24, 14, 13, 23, 27, 30, 46, 12, 7, 13, 32, -18, -2, -10, 1, 18, 6, 6, 32, 19, 11, 18, -10, 30, 41, 37, 33, 9, -6, -26, -32, 9, 31, 0, 29, 39, 1, 46, 22, -1, 14, -20, -12, -3, -5, 67, 36, 56, 53, 33, 17, 69, 35, 13, 39, -8, 4, -22, -19, 3, 29, 35, 51, 31, 30, 36, -1, 1, -3, -13, -5, -8, -6, 46, 82, 74, 77, 74, 72, 43, 31, 7, 9, -3, 11, 22, 15, -10, 42, 42, 64, 58, 72, 26, -20, -13),
  94 => (7, -10, 3, 16, -5, -5, 18, -17, -4, 4, -15, 11, 9, -15, 4, -1, 35, 17, 17, 36, 61, 9, -14, -16, -2, 11, 0, 5, -16, -4, -15, -4, -1, -15, -4, -2, 10, -15, -20, -44, -25, -25, -40, -54, -50, -20, 2, -5, -28, -7, 10, -29, -12, -1, -5, 15, 18, 20, 15, -6, -15, 7, 10, -19, 16, -4, -32, -17, -46, -50, 17, 36, 34, 0, -8, -9, -21, -8, -45, -22, -23, -31, -19, -17, 20, -20, 13, -11, 14, 11, -3, 5, -34, -15, -52, -91, -43, -33, 19, 51, 44, 4, 2, 15, 2, -9, -13, -13, -29, -23, 8, -5, 17, 6, -18, -18, 4, 4, 10, 9, 9, -92, -89, -100, -38, 8, 4, 25, 46, -2, -2, -8, -4, 17, -5, -28, -34, 9, -6, -17, -13, -5, 9, -10, -6, 3, 2, 5, -3, -13, -26, 13, 19, 5, -36, -23, -12, -29, -36, -2, 34, 36, 32, -14, -49, -2, -1, -1, -10, 11, 16, -16, -3, -1, 11, -55, -13, 22, -7, 33, 13, 3, -16, -18, -31, -19, 9, 8, 22, 15, 34, 13, -16, 9, 7, 3, -15, 11, 12, 1, 4, 7, -34, -35, 7, 48, 1, -3, -36, -37, -8, 13, -5, 33, -8, -4, -9, 5, 1, 4, -8, -20, -1, -9, -5, 11, -18, 3, -2, -10, -47, -5, 41, 8, -21, -59, -66, -4, -15, 4, -6, 21, 16, -14, -13, -13, -20, -19, -10, -27, -1, -33, 2, -14, -10, 12, 10, -5, -29, 18, 47, -43, -32, -7, -16, 10, 15, 13, -22, -16, -8, 0, -19, 16, 23, 40, -24, -19, -10, 1, 4, -10, 8, -16, -11, 7, -15, 16, 38, 10, 16, 51, 40, 12, -1, -16, -39, -35, -26, -5, -29, -31, -20, 23, -25, -17, -13, 1, 9, -8, -5, -14, -12, -35, -16, 11, -13, -20, 4, -12, 0, -16, -17, -36, -20, -19, -13, -7, 0, -9, 8, 32, -46, -51, -18, 29, 11, -1, -5, 5, 16, 9, -32, -63, -72, -88, -31, -44, -83, -50, -24, -20, 3, 9, 11, 39, -1, 6, 17, 23, -22, -43, 3, 18, -12, -19, -19, 4, 26, 2, -46, -46, -33, -58, -32, -48, -29, 6, 18, 0, 9, 15, -3, 35, 21, 14, 7, 53, -36, -39, -1, 17, 20, 7, -17, -5, 36, 31, -25, 3, 26, -8, 19, 15, 54, 40, 52, 30, 45, 38, 23, 47, -15, -9, -6, 38, -12, -29, -30, 3, 16, 9, 20, -4, 29, 1, 5, 57, 63, 34, 63, 51, 51, 50, 48, 44, 42, 23, -5, 1, 5, -6, 7, -26, -31, -1, -18, 2, -15, 6, 0, 2, -10, 37, 34, 57, 58, 37, 34, 16, 26, 22, 11, 10, 6, 7, -8, -17, -18, -12, -6, -14, -33, -46, -44, 21, 17, 19, -16, -9, 4, 17, 23, 56, 26, 30, 17, 9, 26, 37, 12, -5, -10, -16, -33, -10, -21, -1, 6, 19, 10, -26, -27, -30, 15, -17, -17, 17, 3, -21, 9, 43, 18, -35, -20, -10, -33, -20, -25, -33, -80, -62, -51, -23, -25, -12, 19, 32, 6, 6, -48, -31, -18, 10, -13, 4, -36, -36, -66, -71, -96, -84, -123, -128, -134, -93, -57, -33, -57, -65, -31, -5, -36, -28, 18, 21, 22, 7, -28, -44, 9, -3, 0, 16, -8, -37, -118, -106, -92, -118, -123, -126, -128, -129, -57, -31, -21, 15, 12, 4, 4, 2, -21, -1, 15, -29, 0, -18, -10, -4, 10, -12, 7, -45, -83, -62, -75, -72, -92, -99, -53, -21, -18, -19, -7, 57, 38, 2, 4, 8, -7, 13, -2, -67, -27, -8, 11, -2, 20, 11, -34, -21, -5, -5, -16, 12, -7, 16, 23, 19, 19, 9, 19, 57, 79, 61, 0, 28, 7, 10, 21, -10, -54, -32, -2, 14, -2, -17, -13, 8, 22, 36, 63, 62, 53, 23, 37, 18, -7, 18, 14, 39, 46, 40, 14, -22, -39, 30, 34, -64, -59, -39, -17, -4, -13, -1, -8, -1, 55, 80, 65, 29, 15, 5, 13, 17, -17, 2, 31, 44, -2, -15, -13, -21, -48, -15, -13, -31, -19, 5, -18, -3, 16, -12, 33, 46, 24, 47, 51, 34, -3, -1, 18, 24, 38, 19, -2, -8, -38, -34, -33, -64, -34, -53, -68, -56, -39, -61, 8, 20, -1, -7, 4, 16, 30, 39, 60, 51, 3, 46, 25, 55, 15, 29, -7, 0, -28, -39, -30, -15, -18, 17, 14, -58, -51, -46, 12, 7, -10, 15, -17, 21, 0, 1, 17, 1, 20, 16, 7, 33, 43, 37, 4, -15, -31, -26, -2, -26, 6, 5, -8, -13, -39, -40),
  95 => (11, -15, -18, 4, -8, -10, 16, 19, 0, 12, 20, 9, 19, 20, -2, -2, -3, -21, -3, 4, -9, 25, 18, -19, -4, 14, 11, 13, -1, 9, 2, 19, 3, 19, 11, -10, -8, -8, -21, 10, 2, -8, 7, -27, -24, -50, -40, 11, 19, 30, 7, -1, -13, -11, 7, -15, -5, -1, 14, 5, 7, 17, -7, 10, -10, 5, 5, -3, -21, 3, -15, -28, -21, -26, -46, 21, 18, 40, -2, 26, -32, 21, -11, -12, 11, -19, -5, -6, -2, -16, 1, -6, 12, -11, 2, 28, 34, 28, -9, -7, -21, -36, -2, 38, 16, -11, -31, 8, -14, -8, 20, -9, 9, -4, -4, -7, -20, -5, -11, -17, 13, 8, 7, 25, 28, 13, 4, -1, 8, 20, 33, 58, 34, -6, -8, 45, 10, -46, -4, 14, 14, -7, 3, -5, -3, -12, 13, -1, -11, 9, 1, -12, -24, -20, -36, -13, 9, 0, 19, 26, 38, 10, 9, 22, 61, -6, 0, -11, -18, -19, 11, 1, 4, 12, 10, -17, 16, -59, -50, 2, -14, -62, -28, 7, 7, 11, 47, 14, -15, -18, 17, 56, -4, -41, -19, -8, 4, 10, 9, -7, -18, 19, 3, 8, -41, -83, -23, -6, -46, -85, -35, -29, 30, 36, 16, 30, -3, 9, 21, -2, -32, -52, 21, 15, -7, -14, -3, -8, -13, 18, 7, -20, -41, -20, 4, -37, -36, -44, -5, -3, 28, 15, 8, 4, 27, 17, 13, 18, -47, -56, 1, 16, 2, 2, 18, 14, 10, -14, -17, -22, -42, 18, 14, -49, -62, -38, -52, -45, 9, 16, 6, 28, 36, 19, -33, -35, -56, -60, -3, -2, -15, 10, 6, -1, -11, 13, -21, -10, 6, -9, 17, -66, -66, -83, -55, -44, -24, 29, 32, 12, 7, 15, 13, -24, -16, -68, -44, -29, 10, -2, 18, -7, 4, 6, -1, -5, -3, 23, 15, -60, -74, -82, -69, -21, 29, 49, 21, 13, -3, -22, -20, 3, -22, -13, -40, -20, -7, -17, 10, 11, 13, 16, -12, -47, -79, -54, -77, -82, -59, -20, -31, -10, 37, -7, 14, 17, 27, 12, 6, 29, -24, -23, 14, -19, 1, -6, 3, 20, 16, 6, -13, -25, -87, -117, -119, -64, -32, -13, -1, 4, 41, 4, 3, 20, 36, 34, 46, 33, -20, 3, -30, -73, -2, -12, -18, -13, 12, 10, -8, -33, -73, -110, -102, -69, -30, -57, -37, -9, 21, 12, 12, 22, 67, 41, 28, -1, -38, -3, -38, -60, -14, 10, -13, -11, -9, -15, 6, -47, -105, -75, -54, -36, -56, -87, -24, 26, 29, 29, 51, 31, 37, 7, 26, -29, -33, -2, 28, -44, 14, -15, -9, -1, -3, 9, -3, -53, -121, -94, -42, -22, -80, -47, -32, 19, 19, 55, 52, 36, -3, 11, -5, -7, -45, -1, 3, 0, 0, 2, 9, -15, -3, 8, -20, -77, -71, -29, -41, -17, -23, -24, 5, 2, 50, 71, 34, 22, -25, 8, -18, -5, -25, -13, -52, -49, 4, -13, 7, 19, 18, -14, -26, -49, -55, -49, -20, 0, -18, -15, 27, 25, 65, 31, 25, -2, -5, 3, -28, -28, -10, 7, -23, -39, -17, -4, 8, -15, 19, -18, -17, -60, -46, -17, 23, 9, -19, 6, 24, 42, 34, 44, 26, -2, -36, -34, -34, -42, -40, -8, -42, -37, -4, -19, 4, 4, -1, -33, -30, -27, -22, -10, -18, 35, 24, 29, 55, 25, 26, -6, -4, -27, -47, -23, -37, -54, -52, -55, -25, -53, -14, 0, -2, 3, -3, -1, -37, -57, 13, 11, -2, 52, 19, -16, 67, 69, 8, 13, 9, 13, 29, 25, 8, -9, -13, -37, -34, -27, 13, 17, -10, 2, -38, -9, -28, -1, 16, -1, -18, 35, 56, 37, 45, 76, 48, 30, 26, 14, 12, 19, 29, 8, -25, -25, 15, 9, -2, 15, -6, 19, -26, 3, 13, 14, 31, 51, 50, 93, 81, 66, 35, 31, 50, 13, 9, 18, 23, 23, -28, -47, -56, -5, 8, -8, -13, -18, 16, -15, 23, 54, 55, 66, 84, 93, 75, 59, 98, 47, 44, 48, 7, 17, 29, 11, 19, 6, -43, -33, -34, 0, 1, 24, -8, -16, 11, 6, 2, 81, 66, 62, 67, 43, 24, 40, 75, 23, 43, 36, 12, -8, 22, 1, -29, -40, -24, -8, 6, 27, 44, 32, 2, 14, 20, 6, 7, 18, 71, 63, 40, 40, 15, 46, 67, 13, 9, 32, 13, -5, -13, -14, -18, -35, -12, -22, 27, 22, 29, 24, -15, -3, 17, -20, 10, -17, -10, 58, 21, 47, 12, 1, 25, 29, 29, 14, -13, -40, 9, 50, -8, 9, -7, -27, 20, 11, 50, 81),
  96 => (-1, 18, 9, -14, 10, 4, 1, 8, -5, 7, -8, 4, 11, 12, 29, -6, -14, 18, 30, 56, 35, 14, -11, 10, 9, 1, 6, -7, -7, -1, 1, 3, 15, -20, -11, 8, 18, 20, 32, 20, 3, 14, 26, -31, -37, -2, 27, 32, 24, 22, 19, 8, -5, 3, -11, 10, 18, 4, -3, 14, -18, -16, 13, -20, -18, 43, 11, -3, 5, -23, -27, -28, 6, -6, -14, -18, -33, -24, 5, 1, 20, -11, 15, 14, -11, -19, -20, 7, -5, 17, -6, 9, 34, -11, -29, -21, -11, -2, -1, -25, -3, -18, -10, -23, -7, -33, -11, -23, 28, 25, 16, 13, -12, -6, 5, -12, 19, 6, 9, 16, 14, 16, 31, 17, 26, 15, -23, -26, -37, -37, 19, 14, 5, -17, 3, -31, -5, 10, -19, -9, 16, -6, 17, 3, 3, 8, 3, -12, 39, 6, -11, -3, -32, -18, 11, 1, -9, 9, -5, -8, 10, 8, 8, -17, 4, -7, 5, -8, -18, -15, -1, -19, 15, -15, -13, -33, 11, -1, -19, -19, -28, -18, 3, 21, 22, 2, 19, -20, -15, 12, 9, -4, 9, -3, 16, -13, -21, 10, 4, 14, -18, 18, -42, 15, -17, -37, 18, -15, 2, 30, -6, -2, 13, 37, 18, 13, -14, -38, -7, -12, 9, -7, 56, -10, 12, 17, 15, 1, -12, -9, -44, 15, -11, 3, -3, 37, 38, 12, 22, 15, -19, -29, 14, 14, 2, -36, -15, -23, 33, 4, 52, -1, -20, 12, 16, -8, 7, 3, -29, -3, -17, -44, -10, -20, 3, 28, 25, 12, -21, 10, -12, -4, -6, -6, -4, -34, 11, 27, 45, 31, 6, 11, -15, 1, 18, -19, -28, -73, -43, -23, 4, 10, -8, 17, 40, 3, -19, -26, -20, -26, -37, 14, 22, -8, -14, 23, 3, 58, -4, 6, -6, 10, -18, -5, -48, -22, -3, 40, 58, 49, -12, 21, -19, -23, -33, -13, -22, -31, -45, -44, -19, -16, -9, 64, 7, 47, 9, 10, -13, -5, 9, -17, -31, 15, 26, 45, 57, 48, -11, 8, 17, -21, -19, 15, -5, 2, -39, -36, -15, -17, -20, 42, 24, -27, -12, 11, -18, 10, 24, 25, 43, 12, 39, 35, 31, 32, -2, -10, 21, -7, 4, -2, -15, -25, -57, -44, -43, -26, 16, 46, 17, -38, -13, -8, 17, -17, 44, 32, 18, 36, 58, 52, -9, -2, -24, -16, -27, -37, -37, -36, -32, -7, -33, -8, -10, 4, 55, 54, 32, 0, 11, -17, -21, 5, 43, 46, 9, 19, 27, 14, -20, -49, -45, -61, -41, -58, -73, -44, -26, -18, 19, -2, 6, 31, 59, 62, 2, -6, -11, -4, 17, 12, 8, -24, 15, -61, -48, -56, -52, -91, -90, -93, -78, -88, -71, -45, -34, -2, 3, 25, 38, 56, 59, 77, 54, 24, -2, -11, 3, -16, 10, -31, -70, -76, -105, -66, -74, -64, -109, -67, -56, -41, -20, 3, -10, 23, 22, 20, 35, 30, 18, 65, 51, 63, -15, 11, -11, -19, -14, -27, -65, -90, -73, -47, -12, -46, -65, -31, 20, 30, 46, 43, 63, 47, 28, 21, 18, 12, -4, 45, 37, 47, -4, 10, -15, -12, -26, 19, -15, -46, -47, -3, -15, -9, 33, 18, 23, 43, 39, 34, 51, 75, 45, -7, -1, -12, -33, 32, 46, 3, 1, 17, 12, -7, -14, 76, 36, 4, 22, 60, 78, 71, 72, 55, 37, 31, 42, 11, 18, 25, 53, 29, -30, -11, -1, 57, 37, 26, 9, 4, -12, 11, 47, 61, 41, 38, 31, 51, 54, 29, 21, 13, 6, 28, 21, 48, 26, 43, 41, -27, 18, 9, 0, 28, 24, 32, -19, -17, 2, 0, 28, 32, 5, -11, 10, 44, 48, 49, 37, 56, 61, 38, 58, 13, 21, 34, 8, -1, -25, 2, -16, 15, 20, 46, -2, 0, 17, -12, 34, 29, -1, -7, 14, 10, 54, 46, 56, 21, -3, -15, 30, 17, 16, -5, -10, -14, -41, -12, -20, -3, -18, 17, -7, -12, 13, -7, 59, 33, 9, -3, 25, 21, 28, 31, 30, 6, -21, -23, -15, -17, -28, -14, -18, -14, 31, 0, -1, -1, -5, 49, 1, 20, 8, 3, 29, 1, 28, 46, 57, 23, 6, 11, 63, 27, 10, 12, 9, -15, -31, -34, -54, -35, -2, -14, -31, 7, 9, 92, -15, -20, -17, 8, 16, -4, -1, 31, 52, 53, -9, 19, 18, -4, -8, -39, -13, -46, -13, -20, -51, -24, 6, 8, -11, 13, 27, 82, 1, -6, -9, -20, -5, -4, -43, -56, -30, 19, 30, 24, 44, 23, -16, -58, -59, -46, -20, -12, 31, 24, 51, 22, 20, 19, 32, 71),
  97 => (-16, -16, 3, 6, 2, 13, -16, 10, -2, 7, -1, 2, -8, 2, -3, -8, 70, 6, -18, -20, -38, 5, 1, -10, 6, -7, -6, 7, 18, 12, 0, -20, 7, 16, -12, -3, 7, 14, 7, 1, -10, -12, 41, 66, 8, 6, 20, -31, -31, 1, -32, 5, -1, -9, -18, 3, 3, 3, -7, -13, -11, -2, 7, -5, 5, 43, -6, -27, 9, 0, 19, 10, -37, 0, -3, -28, -43, 32, 21, 30, 47, -4, -7, 19, -11, -2, -4, -18, -16, 17, -16, -3, 40, -15, -25, -11, -19, 13, -9, 8, 29, 29, 25, 41, 16, 52, 56, 45, 45, 11, -1, 9, -17, -14, -19, -19, 11, -13, 7, 6, 25, 7, -6, -5, 15, -15, 22, 21, 33, 19, 9, 25, 51, 46, 55, 51, 44, 27, -13, 17, 20, -3, 8, 14, -4, 1, -11, 21, -14, 18, 39, 34, 17, 21, -3, -10, 28, 8, -1, 20, 7, 44, 12, 29, -7, -8, -16, -6, 19, 7, -8, 15, 0, 5, -10, -17, -5, 15, 13, 9, -1, -16, -2, -16, 15, 19, 16, 23, 35, 12, 39, -8, -44, -12, -21, -12, -4, 19, -3, -10, -7, 17, -29, -22, -17, -35, -8, -15, -11, -16, -8, -19, -20, 8, -2, -12, -15, -20, -57, -73, -75, -28, 3, 12, 11, 16, 20, -19, 2, 10, -44, -33, -10, -50, -30, -30, -59, -45, -37, -57, -55, -98, -71, -78, -96, -96, -108, -65, -60, -36, 19, -1, 6, -13, -14, -19, 0, -6, -43, -46, -32, -15, -4, -17, -42, -44, -41, -40, -62, -81, -67, -99, -144, -112, -100, -81, -44, -21, -34, -46, 21, 10, 0, 6, -16, -5, 4, 5, 16, 45, 48, 44, 25, -5, 28, -2, 6, 19, 0, 1, -18, -18, -20, -21, -41, 1, -35, 4, 16, -13, 2, 18, -15, 37, -34, 18, 30, 36, 18, 0, 25, 8, 26, 23, 38, 29, 47, 65, 61, 63, 46, 19, 17, 29, -7, 36, 19, -5, -10, -14, 12, 8, -40, 24, 60, 45, 8, 33, 49, 23, 40, 34, 56, 55, 61, 92, 81, 86, 68, 18, 3, 13, 9, 8, 3, 16, 16, 7, -11, -14, 16, 33, 20, 15, 26, 22, 63, 44, 31, 23, 33, 41, 53, 63, 43, 46, 70, 45, 32, -8, 4, -5, -19, 3, -11, 19, 17, 7, 43, 37, -5, -5, -14, 1, 35, -17, -8, -15, -32, -23, -3, 1, -10, -9, -9, -4, 24, 28, 47, -21, 10, -15, 11, -14, 6, 11, 40, 41, 0, -69, -2, 23, -22, -11, -24, -19, -24, -23, -3, -63, -46, -34, -52, -22, -14, 45, 53, -17, -8, -20, 20, 13, -30, 3, -22, 1, 5, 4, 29, 16, -12, 0, -2, -19, -11, -4, -26, -20, -52, -41, -44, -56, -3, 8, 31, -44, 4, 20, 4, 8, 17, -38, -45, -3, -5, -2, 4, 6, 1, 15, -11, 2, 0, 18, 3, -15, -33, -33, -22, -47, -48, -1, 7, -34, 5, -7, 18, -6, 29, -50, -48, 1, -3, -15, 7, 24, -2, 16, -12, -3, -12, -24, 4, -9, 7, -21, -16, -49, -50, -37, -26, -21, -13, 11, -14, -19, -35, -49, -59, -19, -16, 5, 10, 4, 38, 7, 27, 34, 8, -9, -27, -23, -4, 5, 23, -4, -15, -25, -61, -34, -11, 18, -17, 11, -18, -68, -24, 3, -14, 19, -22, -13, -34, -18, -9, 30, 14, 9, -12, -29, -16, 6, 2, 0, -7, -32, -48, -3, -2, 20, -1, 9, 30, -20, -26, 5, -24, -18, -31, -8, -21, -13, -19, -5, -21, -32, -48, -35, -14, -23, -23, -19, -45, -34, -16, 9, -13, -4, -20, 16, -7, -33, -34, -41, 5, -25, 18, 25, 5, 25, -11, 17, -26, -28, -55, -8, 8, -3, -33, -11, -22, -33, -19, -5, -17, 2, -10, -20, 2, -35, -19, -31, -14, -11, 15, -12, -20, -22, -22, -1, -20, -27, -32, 0, -36, 5, 1, -14, -22, -21, -22, -33, -11, -12, -18, -5, -38, -9, -34, -28, -41, -32, -30, -15, -15, -18, -4, 23, 7, -23, 5, -13, -58, -55, -7, -15, -34, -29, -13, -16, 7, 18, 15, 16, -15, -13, -27, -23, -48, -38, 0, 4, -5, -17, -8, 13, 3, -22, 3, -13, -10, -19, -16, -6, -51, -31, -37, -28, 2, -4, -11, 5, 5, -31, -12, -54, -36, -45, -11, -4, -6, -26, -4, -19, -3, -32, -11, -8, -25, 14, -18, -64, -6, -7, -7, -2, 7, 12, 10, -16, 7, -28, 2, -16, -49, -28, -37, -9, -12, -23, 23, -4, 2, -5, -36, -23, -27, 3, -48, -25, -2, 12, -19, -3),
  98 => (-20, -17, 9, -9, -17, -8, -15, 13, 5, 18, -20, 10, -8, -7, 21, 2, -6, 6, -11, -2, -28, 19, -14, -14, -11, -4, -20, -16, -12, 1, 13, 17, 19, -21, 15, 0, -6, -15, 6, 20, 71, 44, 41, 2, 50, 51, 27, 60, 26, 26, 51, -8, 19, 0, 3, -5, -20, 12, 10, 3, -9, -4, 16, 3, -5, 25, 32, 70, 71, 39, 28, 15, 32, 45, 75, 86, 86, 57, 30, 39, -14, -30, -2, 20, 13, -20, 12, -16, 2, -4, -10, 14, 43, 73, 116, 93, 100, 54, 28, 17, 57, 61, 44, 67, 77, 63, 64, -4, -13, -37, 4, -11, -6, 6, -19, -6, 3, 13, -14, 22, 48, 29, 80, 96, 47, 29, 32, 6, 75, 70, 61, 59, 57, 30, 38, 56, 1, 1, -15, -13, 1, -17, 0, -9, -10, 6, 39, 42, 2, 2, 25, 71, 30, 21, 57, 56, 81, 64, 98, 89, 42, 53, 0, 54, 42, 26, -12, 3, 16, 0, 19, -11, 4, -8, 37, 65, 6, 82, 3, 10, 27, 24, 62, 45, 44, 55, 50, 40, 40, 23, 23, 26, -7, -26, -20, 7, -13, 12, -10, 15, -10, -8, 55, 63, 70, 39, -1, 12, 29, 36, 0, 44, 26, 42, 48, -4, 22, 29, 34, -1, 14, -13, 4, -8, -2, 11, 9, -14, -2, 13, 58, 51, 59, 12, -5, 11, -11, -1, 8, 35, 1, 31, 20, -12, 0, -15, -47, -25, -64, -54, -15, 12, 2, -13, 3, -15, -11, -14, 92, 31, 1, -11, 18, -14, 20, 47, 61, 29, 22, 32, 51, 24, -4, -23, -36, -50, -45, -64, -44, -34, -19, -5, -1, -15, 17, -40, 13, 5, 0, -23, 7, 31, 36, 37, 32, 26, 16, -22, -26, 2, -37, -41, -15, -21, -41, -25, -10, -20, -5, 1, 2, 16, -18, -88, -64, -44, -47, -4, 26, 28, 50, 52, 14, -5, -7, -4, -25, -23, -72, -47, -7, -15, -24, -5, -5, 12, -4, -7, -17, 4, 2, -49, 5, -18, -17, 12, 46, 41, 33, 33, 7, -36, -18, -24, -36, -15, -8, -68, -27, -12, -3, -46, -11, 5, 15, 8, 20, -5, -4, -27, 14, -11, -5, 17, 13, 35, 55, 65, 26, 9, 1, -14, -19, -15, -10, -33, -27, -21, 11, -9, -33, -12, 9, -3, -20, -9, 25, -23, 26, 27, 3, -9, 13, 11, 2, 21, -21, -21, -30, -19, 0, -12, 22, -33, -22, 13, 14, -24, 2, -16, -9, 10, 19, 16, -4, -12, 20, -14, 1, -24, -10, 15, 14, 0, -19, -28, -15, -2, -35, -11, 53, 39, 3, -27, 0, 9, 10, -13, -19, -10, 0, -9, -42, 8, -15, 28, -16, 17, 10, 11, 33, -2, -24, 2, 0, 21, 9, 12, 29, 34, -4, -30, 5, 45, 33, -9, 11, -14, -5, -3, -6, 2, 14, 57, -18, -13, 23, 10, 22, 16, 9, 21, 12, 21, -15, -3, 35, 52, 36, 3, -7, -1, 34, 2, -16, -3, 5, 15, 38, -22, 4, 11, -15, -1, 24, 18, 14, 58, 21, 39, 3, 16, 6, -14, 10, 40, 30, 27, 21, -7, 47, -32, -16, -6, -15, 18, 11, -29, 25, 5, 4, 11, 19, -11, 16, 28, 18, 23, 38, 47, 11, 9, 8, -1, 39, 6, -17, -5, 29, -29, -15, -6, 20, -9, 50, -17, 30, 39, 4, -4, 27, 10, -12, 13, 14, 13, 40, 11, 19, 43, 15, 31, 44, 46, 45, 24, 12, -41, -9, -3, 18, -13, 38, 47, 101, 55, 2, -11, 19, 44, 29, 47, 59, 59, 44, 57, 45, 64, 77, 68, 71, 59, 56, 28, 35, 27, 10, -18, 6, 10, 34, 25, 54, 85, 12, -10, -1, 41, 53, 55, 37, 47, 70, 88, 36, 61, 54, 48, 69, 61, 53, 53, 61, 55, -8, -14, -10, -19, 48, 31, 62, 60, 62, 52, 37, 25, 69, 48, 47, 20, 52, 28, 46, 36, 36, 33, 44, 31, 42, 64, 25, 60, 16, 19, 6, 6, 17, 2, 10, 49, 44, 62, 52, 43, 28, 50, 41, 23, 50, 63, 32, 47, 46, 57, 29, 27, 38, 21, 21, 13, -1, -10, 12, -1, 3, -18, 18, -10, 19, 31, 43, 16, 20, 49, 36, 40, 64, 18, 27, 29, 23, 29, 19, 23, 10, 12, 1, 28, -13, 11, 6, 19, 6, 10, -24, 4, -7, -9, 6, -17, 27, -3, 15, 1, -12, -28, 8, -21, -10, 4, 30, 44, 5, 14, -14, 18, -1, 15, 15, 13, -10, 25, 5, 44, 44, 31, -11, -16, 23, 45, 9, 33, 22, 33, 26, 47, 26, 37, 79, 56, 58, 14, 31, 15),
  99 => (-11, -3, 1, 8, 5, 9, 1, 13, -16, -13, -7, 3, -16, -3, 53, 46, 30, -22, -2, -6, -20, -30, 11, 18, -10, 15, 9, -12, 19, 20, -13, 11, -8, -19, 10, 14, 10, 9, -19, 8, -8, 51, 15, 24, 43, 1, -4, 16, 35, 10, 33, -36, 20, -12, -3, -20, 9, -20, -7, 2, 7, 4, 14, 2, 15, -22, -28, 1, 9, 30, 37, -5, 11, -19, -6, -2, -18, -15, 4, -2, 24, -9, -10, -13, 6, -18, 10, 16, 0, -20, 17, 18, -3, -15, 0, 53, 64, 7, 3, 10, 15, 10, -21, 13, -20, -57, 2, -26, 2, -14, 0, 14, 16, -18, 5, -6, -8, 18, -15, -9, -23, 43, 62, 41, 10, 6, 15, 27, 40, -4, -10, 16, -17, -27, -14, 4, -25, -22, 20, 11, 0, 15, 5, 3, -10, -5, 1, 10, 10, 33, 38, 25, 17, 8, -22, 58, 22, 13, -28, -13, 15, 11, 3, -10, 31, 0, 5, -5, -2, 10, -11, -18, -14, -3, 10, -1, 25, 33, 24, -14, 30, 10, 0, 22, 27, 10, -2, 8, 7, 30, 16, 29, 40, -6, -24, -15, 18, -1, -2, 4, 18, 3, 11, -1, 5, 27, -1, -22, 20, -37, 4, 23, -19, 13, -16, -2, -6, 19, 21, -1, 18, 9, -41, 18, 10, 7, 19, -15, 6, -11, 39, 27, -4, 23, 23, 23, -25, -37, -26, -10, -13, -6, 25, 32, 19, 14, -8, 19, -1, 13, -19, 0, -6, 20, 12, 10, 12, -2, 16, 4, 18, 32, 13, 32, -8, 23, 27, 13, -26, -15, 36, 25, 43, 1, -16, 11, 41, -10, 12, 31, -11, 18, 5, -18, 11, 24, 13, 5, 4, 53, 59, 64, 47, 36, 40, -11, -23, -33, 24, 4, 45, 6, 13, 5, 40, 1, 37, 27, 2, -6, 5, 20, 13, 30, 0, -27, -14, 58, 56, 48, 47, 10, 29, -15, -41, -10, 14, 11, 35, 51, 41, 15, 13, 9, 23, 32, -12, 18, 0, 8, 13, 6, -16, -33, -12, 32, 74, 51, 44, 20, -7, -48, -79, -12, 7, 17, 35, 15, 13, 16, 17, 42, -23, 43, -12, 6, -19, 15, 17, 9, -44, 2, -12, 62, 62, 40, 9, -35, -11, -4, -36, -24, 27, 25, 42, 40, -25, -27, -3, 17, -62, -10, -18, -14, -10, -18, -2, 31, -3, 2, -23, -1, -15, 10, -55, -85, -58, -59, -92, -70, 0, 13, 7, 8, -19, -42, -3, 32, -38, 15, 8, -14, 0, 10, 22, 19, 35, -11, -33, -72, -126, -118, -95, -98, -81, -106, -97, -42, 15, 17, 4, -20, -27, -42, -9, 20, -46, 35, 10, -15, -3, 0, 28, 39, 2, 9, -22, -41, -94, -61, -25, -48, -67, -70, -54, -34, -9, -21, 0, -8, -1, 11, -16, 37, -5, 16, -5, -4, 3, 16, -11, 30, 3, 9, -23, -15, -52, -60, -68, -38, -67, -87, -82, -28, -11, -19, -2, 18, -6, -6, -24, -13, -31, 20, 15, -1, -10, 10, -12, 35, 31, 33, 2, 11, -71, -62, -88, -34, -42, -46, -46, -14, -5, 20, 32, 11, 21, 1, 17, -17, -27, 59, -19, -9, 9, -6, 24, 3, -5, 20, 33, -21, -29, -35, -64, -81, -91, -40, -5, -4, -31, -21, 10, -7, 31, 6, 9, -9, -2, 72, -2, -12, -14, -15, 0, -10, 8, 34, -3, -35, -56, -38, -23, -63, -64, -34, -42, 9, 14, 17, 16, 11, -19, 13, 3, -6, -30, 80, -19, -11, 18, 4, 2, -37, 16, 18, 20, -44, -24, -39, -64, -19, 11, 27, 11, 30, 1, 28, 32, 13, 17, -11, -18, 0, 10, 57, 10, 1, -14, 5, -16, -15, 15, 8, -7, -23, 12, -6, -19, -27, 5, 8, 15, 31, -1, 9, 23, 54, 40, 29, 4, -30, -4, 48, -18, 14, -13, 0, 3, -10, 22, 18, -2, 5, 17, 51, 58, 28, 26, 27, 13, 43, 35, -9, 43, 26, 63, 10, 20, -41, -13, 72, -7, 3, -2, 1, -41, -34, -12, -11, -11, -15, 5, 43, 72, 39, 61, 40, 24, 18, -12, 14, 53, 28, 31, -9, -4, -10, -12, 56, 0, 5, -8, -13, 2, -51, -30, -21, -8, -31, -26, -28, 20, 18, 35, 43, 25, 11, 33, 43, 53, 51, 9, 3, 22, -9, -17, 46, -20, 14, 18, -1, 18, -21, -8, -9, -6, -20, -38, -44, 19, 43, 35, 43, 26, 24, 28, 63, 71, 52, 71, 12, 3, -7, 19, 0, 3, -7, 5, -9, -18, 18, -9, -18, -18, -13, -22, -29, -22, -6, 6, 26, 6, -3, -15, 11, 21, 55, 75, 52, 1, -11, 20, 5),
  100 => (-9, 14, 1, -3, -20, -15, 4, 0, 15, 10, 1, 15, 5, -15, -1, 31, -35, -7, 19, 33, 23, 17, 23, 8, -15, -1, -12, 8, 8, -3, 2, 6, 8, 9, 0, 9, 16, -7, -15, 7, -8, 25, -5, 40, 59, 67, 14, 17, 51, 5, -3, -15, 6, -18, -16, -16, 19, 15, -10, 14, -12, 6, 8, 11, 17, 4, -15, -21, -32, 27, 36, 7, -3, -21, -2, 0, -16, 19, -17, -20, -13, 2, 2, 3, 3, -8, -4, 12, 15, -5, 7, -20, -2, -6, -18, 3, 3, 1, -20, 14, 6, 14, 9, -3, -4, -13, 8, -6, 13, 24, 10, -18, -8, 20, 2, 1, 1, -14, -15, -35, -29, -41, -63, -36, -12, -83, -53, -14, 12, -12, 22, -26, -11, 1, 20, -3, -16, 4, 12, 12, 8, -9, -4, -15, -20, 19, -42, 10, -33, -23, -10, -10, -6, -96, -35, 14, 39, 23, 21, -37, -9, 0, 3, -33, -53, -9, 9, 12, -15, -17, -4, 4, 2, 11, -9, -33, -33, -28, 14, 32, -22, -55, -16, 40, 38, 14, 24, -19, -4, -3, 9, -29, -21, -39, 26, -13, -1, -20, -19, 8, 18, -18, 4, -43, -6, 24, -3, 16, -25, -53, -15, -1, 19, 20, 22, -6, -50, 33, 46, 3, -30, -16, 39, 17, 10, 6, -13, 2, -7, -14, -8, -11, 5, 24, 65, 22, -35, -69, -23, -15, 20, 43, 14, 6, -48, 10, 65, 28, -11, 29, 38, 18, -10, 13, 6, 8, -1, 2, 25, 4, 11, 44, 23, 40, 4, -13, -37, -20, 38, 6, 16, -19, -49, 24, 30, 27, -9, 1, 0, 11, 16, 13, -4, 12, -10, 7, 32, -21, 56, 40, -7, 32, 37, -10, -29, -12, 59, 16, 26, 20, -61, 3, 23, 7, 4, -15, -1, 16, -12, 20, -11, -3, 12, 35, 34, 27, 73, 48, 11, 41, 37, 4, 1, -11, 11, 4, -1, -8, -70, 15, 32, 32, -39, -46, -9, 52, -15, 19, -17, -11, -34, 16, 5, 4, 18, -5, 28, 65, 10, 14, -17, -5, 16, -17, 31, -8, -48, 6, 35, 46, -13, -26, -10, 63, -14, -5, -14, 3, -6, 17, 10, -5, -8, -17, 8, 53, -13, -67, -40, -15, 11, 20, 28, 7, -53, -21, 21, 47, 15, -41, -40, 18, -2, -20, 0, 7, -3, 15, -23, -30, -21, -48, -26, 22, -3, -89, -29, -14, -14, 35, 24, 27, -33, -47, -17, 19, -24, -19, -28, 11, -3, -18, 6, -5, 10, 44, -14, -24, -11, -45, -16, -4, -32, -60, -43, 10, -12, 12, 13, 0, -35, -73, -2, 2, -17, -33, -61, -44, -2, 10, 18, 16, 9, 13, -24, 10, -11, -16, -33, 2, -70, -90, -53, -40, -41, -5, -1, -8, -15, -80, -29, -26, -2, 22, -49, -26, -15, 1, 11, 20, -39, -50, -49, 2, -2, -43, -20, -13, -86, -81, -53, -16, -15, -26, -23, 11, -23, -89, -36, -15, 26, 1, -12, -27, -7, 20, -8, 7, -21, -43, -25, 8, -3, -8, 10, 16, -57, -65, -67, -43, -31, -10, -15, 36, 7, -77, -69, -7, 12, -12, -39, 10, 3, 12, 3, 10, -41, -31, -19, 10, 28, -7, -9, 13, -11, -54, -79, -57, -29, -24, -3, 16, 1, -51, -33, -19, 31, 20, 20, -13, 14, 20, 18, -16, -42, -50, -48, 32, 54, 25, 26, 10, -1, -61, -93, -35, -26, -13, 6, 11, -20, -72, -42, 6, 25, 24, 41, -35, 12, 19, -12, 17, -30, -45, -28, 23, 44, 21, 16, -15, -4, -39, -60, -41, -44, -53, -19, 13, -21, -38, -34, 3, 29, 31, 39, -4, 4, -7, -14, 7, -28, -39, -55, -21, 31, 1, 15, 16, -7, -50, -56, -42, -30, -24, 9, -8, -18, -29, -22, -29, 20, 47, 45, -14, 12, -13, 18, 14, -37, -39, -69, -3, 40, 32, 20, 9, -6, -21, -25, -37, -23, -21, -23, 41, 50, -4, -56, 1, 12, 41, 25, -1, 6, -16, -11, -13, -33, 7, -45, -29, 35, 21, -8, -14, 19, 0, -24, -21, -44, -10, -2, 50, 82, 56, -14, -5, 14, 35, -1, -11, 6, -9, -2, 19, -13, -11, 7, -26, 3, 11, -22, -26, 10, 2, -31, -40, -51, -7, -2, 34, 53, -3, -31, 7, 32, 5, -9, -48, 3, 19, -14, -8, 6, 6, -7, -11, -12, -6, -5, -31, -19, -8, 4, -14, -11, 14, -21, 21, 41, -29, -34, -3, 12, -8, -2, -47, 17, 16, 9, -7, 6, 4, -7, -4, -20, 1, -57, -20, 7, 9, -2, 8, 27, 23, 11, 12, 42, 16, 0, 27, 23, -1, -7, -23),
  101 => (-3, 8, -5, 18, 18, 14, 20, -18, 11, 17, 18, 17, -8, 4, 7, 1, -30, -20, 38, 17, 15, -9, 8, -3, -14, 13, 16, -13, 12, -9, 16, -3, -2, 13, -2, 7, -7, -20, 4, 51, -8, 34, -30, 3, 22, 18, 40, -12, -3, 34, 22, 54, 29, 5, 1, 1, -1, 17, -13, 3, -4, -9, 10, 17, 5, -2, 63, -22, -45, 2, 27, 16, -5, -9, 1, -23, 29, 31, 70, 23, 44, -20, 17, -19, 0, 19, -16, 14, 18, 11, 14, 18, -24, 29, 27, 6, 39, 28, 8, -1, -13, -15, -33, 0, 9, 8, 8, 24, 20, -9, -15, -6, -5, -5, 9, 5, 10, -7, -6, 5, -5, 20, 31, 45, 39, -9, -8, 9, 8, 17, -20, -25, 10, -3, 4, -18, 10, -26, -2, -7, -4, -9, 2, 15, -13, 11, -16, -15, -41, -3, 18, 1, 13, -21, -9, 24, 32, -3, -22, -6, -15, 26, 12, -23, -58, 31, -6, -3, -3, -8, 3, 3, 11, 11, 2, 4, -32, -24, -33, 11, 21, -5, -25, -1, 38, 6, 21, -2, 4, 3, 21, 16, -10, 7, -3, -4, -4, 18, 9, -13, -6, 2, -38, 32, 17, 1, -18, -13, -13, -10, 20, 23, 5, 24, 17, 12, 1, 42, 18, 15, 8, 3, 6, -1, -18, -13, 19, 6, 7, 12, 10, 30, 8, -5, 5, 4, -13, -27, -26, 0, 7, -12, -16, -4, -14, 6, -4, 25, 21, 23, -24, 11, 9, -15, 10, 1, 4, 4, -21, -4, 10, -11, 16, 31, 2, -41, -37, -18, 5, -14, -8, 13, -18, -40, 15, 41, 40, 32, -25, -4, 3, 14, 13, 4, -10, 6, 2, -8, 11, 21, 30, 34, 12, -69, -58, -1, -1, 1, -12, 24, 24, 11, -3, 1, 12, 29, -6, 16, 2, 12, 5, 10, -6, -48, -8, -71, -2, 0, 14, 19, -20, -81, -64, -2, 5, 19, 24, 48, 15, -19, -40, -35, 22, 34, 18, -6, 10, 15, 3, 3, 2, -2, -40, -19, 10, 3, 23, 26, -27, -86, -73, -22, 31, 23, 28, 2, 4, -13, -54, -66, -12, 26, 18, 8, 18, -2, -6, 18, -32, -29, -55, -6, 28, 12, 31, 45, -47, -57, -71, 20, 40, 2, 28, 15, -5, -32, -74, -64, -15, -8, 10, 11, 16, 5, 6, 12, -10, -36, -54, 47, 34, 8, 22, 21, -83, -62, -93, 28, 35, 7, 24, -3, -7, -59, -42, -78, -16, -23, -5, 2, -8, 11, 19, 3, -31, -26, -16, 40, 40, 5, -2, 6, -97, -81, -78, 39, 21, 37, 54, -15, -38, -46, -40, -62, -17, -32, 5, 3, -3, 20, 20, -3, -54, -15, -7, 30, 15, 46, 23, -1, -66, -85, -48, 32, 19, 56, 63, 5, -52, -79, -65, -50, 3, -11, -37, 11, -20, -19, 12, -13, -35, -18, 13, 18, 37, 27, 13, 0, -58, -93, -38, 29, 30, 37, 64, -9, -41, -20, -56, -59, -11, 6, -36, -8, 11, -7, 11, 11, -50, -13, 21, 14, 21, 6, -6, -51, -75, -86, 3, 36, 15, 31, 54, 7, -30, -16, -18, -26, -17, -10, -20, -16, 5, -14, 11, 16, -33, -6, 40, 18, 18, -25, 10, -70, -70, -70, 13, 9, 17, 21, 43, -7, -20, -37, -19, 21, 32, 5, -2, 16, -16, -15, -1, 0, -27, 6, 28, 5, 14, 1, -1, -31, -24, -22, -14, 28, -1, 18, 21, -9, -39, -49, -36, -27, 0, 13, -26, 11, 6, -18, 19, 0, -1, 30, 24, 12, 25, -1, -8, -32, -60, -25, 40, 8, 28, 12, 25, -57, -48, -64, -10, -42, -16, -40, -44, -11, -18, 3, 8, 10, 12, 63, 21, 7, 31, -33, -31, -56, -44, 3, 35, 22, 34, 28, 30, -58, -58, -35, -14, -8, -35, -39, -36, -12, -17, 19, -6, 1, 36, 24, -5, 7, -9, -25, -38, -52, -46, 17, 24, 30, -1, 12, 13, -40, -103, -51, -50, -46, -3, -51, -18, 9, 15, 9, -5, -14, -5, -2, 24, 23, -11, -20, -39, -17, -32, 48, 36, 30, 21, 25, -11, -30, -61, -49, -51, -19, -13, -13, -33, -1, -7, 9, -9, 17, 3, 8, 6, -14, -24, -24, -41, -15, -8, 35, 52, 16, 13, 8, 10, -33, -45, -39, -39, -40, -7, -38, -28, 12, -18, 5, -15, -9, -17, -4, -19, -14, 5, -4, -16, -36, -17, 13, 34, 44, 40, 43, 43, -9, -16, -25, -24, -44, -15, -9, 12, 19, 17, 6, 16, -8, 8, 3, -32, 5, -12, -3, -4, -7, -49, -2, -1, 19, 68, 14, 9, 25, 23, -16, 15, -18, -41, 12, 24, -1),
  102 => (-7, -20, 17, 4, 2, 16, 15, -18, 7, -18, 7, -4, -10, -18, 21, 2, -10, 15, 32, 22, 16, -22, 0, 5, -17, 14, -9, 9, -13, -6, -18, -11, -3, -10, -15, 5, 13, 17, 11, -7, 6, -4, -29, -21, -56, -45, -22, -28, 19, -32, -21, 0, 0, -9, -16, -12, 5, 1, 9, -2, -2, 13, 5, -8, 5, 27, -30, -57, -20, -1, -3, 27, 18, 15, 69, 42, 0, -26, -61, -43, -20, 3, -13, -6, -3, 2, 9, 6, -20, -7, -12, 19, 2, -35, -45, -36, 13, 4, 31, 13, 4, 0, 41, 35, 21, -5, -68, -30, -73, 4, -18, 6, -5, 9, 4, 1, 12, 19, -1, -1, 6, 5, -20, -22, 21, 19, 15, 25, -12, 17, 35, 64, 99, 64, 8, -8, -38, -6, -11, 4, -3, -4, 20, -17, 7, 7, 2, -2, -5, 10, 7, 45, 16, 54, 53, 1, -4, 22, -2, 50, 87, 32, 0, -23, 38, -33, -13, -2, -16, -17, 5, 5, 3, -1, 4, 35, -13, -22, 29, 47, 14, 28, 34, -4, -12, 1, -36, 7, 46, 57, -2, 6, 52, 1, 16, -8, -5, 0, -13, -10, -11, -20, -18, 9, -16, -31, 2, 18, -10, -15, -24, -28, -6, -15, -67, -19, 19, 27, -8, 1, 47, 28, -6, -39, -6, -2, 19, -16, 15, 19, 38, 8, -30, -13, -46, -20, -13, -36, 23, -1, -14, -42, -74, -56, 3, -11, -31, -16, 21, 39, -29, -68, -15, 10, 7, 14, -14, -10, 40, -17, -67, -50, -39, -27, -19, -9, 1, 37, 14, -18, -77, -49, -27, -31, -1, -17, 9, -5, -37, -60, -17, -4, -8, -5, 20, -18, -1, -22, -19, -47, -68, -26, -39, 0, 14, 34, 32, -10, -81, -70, -40, -62, -18, -7, 5, -39, -27, -45, -16, 17, -12, -19, 2, -3, -6, -40, -42, -36, -61, -8, -9, 3, 29, 20, -4, 1, -40, -21, -21, -45, -16, 6, -6, -11, -25, -16, 12, 6, -5, 4, -16, -26, -20, -35, 13, -3, 3, -10, 3, 7, 17, 47, -4, 12, -31, -5, 2, -58, -25, -11, -39, 7, -20, -39, 0, -8, -9, 13, -9, -4, -15, -16, 46, 5, 24, 24, 7, 33, 16, 12, -14, -28, 4, 7, 12, -71, -82, -21, -28, 25, -8, -35, 16, -9, -2, 18, -5, -52, -10, 36, 5, 41, 25, 21, 34, -1, -5, 10, -1, -11, 2, 27, 27, -11, -57, -19, 21, 14, 17, -10, -9, -17, 19, 9, -18, -40, 11, 26, 35, 46, 47, 83, 36, 27, 18, 12, 24, 14, -32, 5, 33, 10, -27, -33, 7, 5, 3, -10, 1, 11, -19, 5, -13, -40, -12, -4, -14, 32, 45, 36, 39, 8, -34, -51, 11, 20, 0, 44, 48, 6, 7, -8, 7, -31, -21, -40, 13, 17, 15, -18, -15, -2, 0, -8, -23, -11, 3, 55, 8, -25, -46, -70, -27, -14, -17, -1, 0, -20, -1, 0, -15, -12, -7, -18, -6, -11, -8, -10, -14, 0, -9, 19, 7, 5, -10, 3, -39, -48, -74, -117, -101, -44, -17, 18, 8, -12, 22, 11, -8, -24, -42, -34, -7, -6, 2, 7, -40, -7, -32, -10, 21, 16, 7, 5, -18, -58, -103, -109, -117, -57, -6, 8, 10, 47, 57, 13, -32, -32, -46, -33, -4, -7, -17, -9, -28, -28, -31, -12, -9, 16, 32, 28, -32, -42, -70, -52, -70, -45, -1, 17, 9, 11, 37, 8, -58, -59, -13, -29, 19, 17, 4, 15, 22, -4, -21, -18, -11, 17, 14, -32, -12, 22, -26, -29, -28, -62, -30, -11, 7, -2, 21, -42, -44, -35, 14, -17, -15, -3, 20, 0, 62, 10, -9, -19, -56, 1, -1, 1, -7, 34, 2, 20, -14, 4, -17, -5, 15, 33, -4, 3, -42, -58, -23, -4, -16, -16, -16, -4, 66, 28, -6, -22, -43, -3, 13, -13, 21, 36, 34, 77, 96, 28, 52, 65, 55, 26, -2, -39, -23, -22, -19, 4, -7, -4, -13, 18, 38, 23, -7, -44, -37, -2, -1, -6, 2, 14, 34, 77, 71, 51, 39, 44, 55, 13, -9, -21, -11, 9, -17, -23, -17, -20, 16, -16, -5, 13, -7, -23, -3, -27, -6, 0, -30, -15, 22, 58, 41, 51, 39, 39, 26, 6, 7, -18, -51, -17, 9, -15, 5, -10, 17, -13, 29, 18, -29, -28, 1, -15, -21, 4, 10, 32, 31, 18, 42, 27, 45, 41, 12, -15, 3, 4, 16, 13, -5, -17, -11, 9, 17, 12, 20, -22, -38, -28, -14, -15, -15, -3, 5, 29, 27, 10, 0, 29, -12, -7, -40, -34, 12, -1, 0, 25, 29, -42),
  103 => (18, -12, 0, 1, -5, 9, 17, -18, 18, 6, 18, -5, 3, -2, 11, 0, -27, -5, 17, -4, -7, 4, 14, -7, -3, -18, -4, 9, -11, 5, -13, -19, 4, -2, 13, -8, -17, -2, 3, -2, -13, -5, -22, 6, 10, 14, 28, 28, -20, -30, -23, 15, 12, -18, 12, -1, -3, -20, 21, -19, 2, 19, 5, 9, -9, 27, 11, -20, 17, -21, -28, -31, -3, 6, -33, -47, -24, -37, 29, -13, 2, -11, 11, -8, 4, -2, -14, 7, 10, -7, 11, 16, 5, -16, -29, 13, -2, -6, -45, -21, -18, -15, -31, -8, -36, -32, 17, 20, -25, -14, -10, 8, 20, 8, 2, -17, -9, 4, -16, 30, 6, -8, -8, -13, -63, -29, -24, 12, -3, -2, -4, -4, 12, 21, 16, -9, 2, -16, -3, 2, 0, 3, 12, 10, 1, -13, 15, -12, -6, -30, -30, -37, -23, -1, 13, 7, -7, -7, 23, 39, 11, 6, 44, -10, -6, 2, 15, -19, 14, 15, -3, 6, -16, 20, -5, 11, 2, -43, 28, 28, 3, 32, 26, 20, 13, 20, 14, 44, 29, 0, 15, 1, 8, -14, -10, -3, -14, -12, -9, 11, 10, -2, -18, 10, 8, -19, 10, 49, 47, 11, 5, 20, 25, -6, 11, -1, -14, -8, -13, -6, 0, -49, -27, 8, 15, 11, -18, 19, -20, -19, 2, 13, 17, -2, -12, -19, -30, -18, -18, -11, 23, -44, -41, -16, 9, -9, -26, -20, -2, -34, -30, -1, -9, -12, 2, -8, -11, 20, -22, 19, -20, 5, -10, -19, -46, -15, -7, -13, 9, 13, -8, -16, -4, -8, -20, -33, 1, -64, -20, 0, 7, -9, 11, 10, -18, -14, -9, 7, 16, 9, 13, 3, -5, 10, 1, -30, -4, 16, 6, -10, 23, 10, -17, 4, -22, -37, -28, -3, -13, 14, -9, -15, 4, 17, -21, -15, 18, 18, -20, -2, 12, 8, -8, -24, 0, 43, 18, -12, -30, -15, -25, -20, -5, -33, -26, 18, -5, -14, 9, -14, 28, 4, 8, -17, -9, -13, -30, -22, -31, -12, -1, 27, 44, 51, 20, 5, -22, -15, -33, -18, 17, 8, 6, 22, 13, 16, 4, 7, 25, -14, -31, -55, -2, -20, -39, -37, -38, -66, -51, -102, -24, -13, -24, 3, 10, -17, 28, 4, 54, 49, 34, -6, -17, -9, 4, -16, 22, 14, -19, -8, -6, 10, 2, -9, -45, -50, -106, -110, -115, -141, -138, -25, -22, -18, -8, 41, 57, 92, 52, 22, 0, 0, 20, 20, 4, 40, 29, 11, 25, 36, 55, 57, 7, 17, -33, -64, -82, -138, -150, -94, -78, -19, 21, 29, 45, 62, 61, -23, -3, -20, -7, 0, 31, 59, -19, 1, -15, -10, 28, 18, 35, 19, 21, -4, -27, -44, -24, -33, -41, 37, 37, -6, 27, 30, 44, -33, -16, 4, -12, -14, 11, 5, -3, -7, -29, -26, -10, 24, -13, 11, -15, 11, 66, 47, 79, 26, 11, 3, 9, 9, -12, 9, 1, -48, 4, 6, -9, 15, 10, -45, 6, -21, -54, -40, -22, -26, -26, 13, 70, 40, 25, 7, 26, 15, -7, -25, -9, -2, -30, -6, 4, -42, -10, 12, 6, 14, 7, -19, -46, -33, -59, -50, -22, -35, -15, -5, 32, 33, 17, 25, 15, -15, 5, -17, 3, -14, -19, -34, -7, -29, 17, 19, 2, -3, -20, -25, -16, -42, -19, -19, -19, -5, -17, -12, 4, 6, 22, 20, 13, 22, 25, -3, -9, -22, -21, -57, -24, -14, 18, 9, 6, -9, 17, 8, -17, -12, 44, 20, 38, 57, 7, 19, 23, 19, -4, 24, 8, 10, 31, 6, 1, 11, -12, -46, -65, -30, -11, 11, 5, 17, 4, 8, 45, 24, 18, 25, 22, 32, 29, 8, 43, 34, 20, -12, -37, 21, 7, -15, -2, 5, -16, -46, -62, -52, 13, 2, -15, -12, -33, 14, 0, 28, 49, 1, 13, 14, 35, 42, 15, 4, 27, 4, -22, 24, -1, -6, -10, 3, -14, -34, -42, -29, -16, -19, -18, -2, -24, 23, 13, 49, 32, 8, 25, -10, 40, 12, -12, -8, 8, -11, 23, 37, -7, 21, -21, 1, 18, -4, -26, -24, -19, 16, 14, 16, -18, 13, -31, -18, 26, 42, -7, 5, 14, 28, 7, 13, 48, 9, 37, 43, -3, -4, 40, -8, 0, -17, -34, -59, 6, 18, 11, -16, -25, -1, -20, -50, -27, -37, -23, 3, 1, -12, 27, 26, 49, 41, 28, 43, 22, 4, -7, -6, -32, -22, -43, -30, 21, -16, -6, -11, 2, -5, -11, -5, -1, -16, -30, -11, -13, -27, -14, -11, -13, -22, 5, -11, 21, -2, 0, 30, -26, -19, -14, -3),
  104 => (-19, 11, 5, -15, 8, 1, 17, 17, 6, 16, 1, -6, -18, 15, 15, -17, -24, -55, -42, -6, 2, 39, -20, 7, 15, 2, -17, -6, -5, -4, -9, -10, -17, -20, 18, 12, -12, 9, 32, 17, 38, 69, 45, 13, 28, -17, -8, 14, 28, 29, 30, 17, 9, 10, 9, -5, -13, 1, 16, -12, 12, -14, 13, 0, 16, -1, 23, 55, 33, 31, -17, -42, -7, 32, 9, -12, -11, 22, 68, 16, 47, 25, -6, 8, 6, 18, -9, 3, -10, 4, -4, -16, 19, 3, -6, -25, -20, -45, -68, -28, 31, 41, 18, 38, -6, 18, 37, -1, 30, 45, -20, -16, -15, 6, 11, 4, -15, 13, 14, 4, 8, 47, 47, 45, 1, -53, -35, -20, 4, 34, -25, 29, 14, 54, 18, 3, 16, 24, -5, 19, -20, -5, -2, 10, -18, -3, 18, 16, 36, 53, 56, 16, -62, -34, -37, -18, -6, 13, -3, -5, 0, 38, -8, -12, -4, 11, 7, 10, -8, -18, 17, -3, 19, 7, -7, 25, 38, 32, 6, 5, -16, -4, -2, 3, -11, 13, -5, -7, 15, 8, 2, 0, 47, -5, 16, -20, -15, -20, -20, -7, -19, -15, 11, 20, 56, 13, 30, 32, -4, -11, 35, 32, 28, 16, 29, -3, 18, 15, 14, -12, 14, 52, 33, 2, -12, 5, -20, 12, 11, 0, 37, 68, 87, 69, 73, 39, 37, -20, 10, 24, 32, 30, 20, 9, 18, 8, 10, 1, 18, 74, 12, -9, 19, 0, 8, 6, 13, -2, 100, 87, 106, 98, 118, 65, 31, -26, -53, 3, -6, 0, -5, 9, 24, 30, 27, 14, 62, 61, 31, 18, -15, 19, 8, -15, 18, 20, 105, 48, 69, 80, 81, 80, 47, -10, -19, 10, 5, -14, 12, 13, 16, 25, 33, 5, 73, 57, 84, 88, -10, 3, 1, -20, -12, 49, 53, 45, 70, 45, 55, 58, 53, 10, -28, -14, 48, 68, 33, 38, 50, 63, 36, 29, 48, 34, 15, 62, -4, -19, 19, 13, -34, -20, -24, 14, 13, -13, 7, 6, 27, 7, -32, -14, -3, -4, -4, 3, -1, -5, 16, 0, 21, -7, -10, 31, -11, -11, -12, -18, -41, -15, -70, -33, 9, 29, 19, 26, 24, 4, 17, -30, -36, -56, -33, -68, -70, -50, -35, -46, -22, -31, 17, -6, 10, 16, 20, -16, -26, -36, -43, -91, -29, -17, -16, 39, -19, -14, -18, -52, -43, -23, -76, -91, -90, -57, -34, -55, -19, 0, 1, 26, -4, 20, -12, 9, -8, -67, -67, -68, -48, -57, -24, -13, -30, -20, -33, -36, 6, 16, -31, -62, -33, -70, -49, -15, -50, -8, -27, -4, -8, 20, 7, 5, -43, -46, -60, -74, -47, -78, -26, -36, -41, -30, -21, -2, -9, 7, -1, 14, -12, -20, -11, 18, 2, 20, -30, 5, -14, -6, 11, -2, -67, -33, -50, -78, -60, -66, -44, -86, -16, -26, -22, -17, -25, 6, -14, 1, -31, -9, -10, 21, -14, -15, 13, 21, -3, -7, -18, 1, -27, -10, -46, -40, -46, -17, -28, -65, -26, -54, 0, -15, -4, 9, 1, 3, 16, -13, -33, -24, -26, -6, 14, 18, 7, 16, -6, 12, 17, 2, -25, 7, -12, -16, -31, -64, -42, -52, -14, -15, -27, -19, -36, -3, -6, -26, -42, -36, -25, -10, -50, 13, 11, 20, -10, -11, 37, -8, -15, 21, 19, 20, 5, 7, 20, -21, 5, 0, 29, 14, -2, 36, 2, -6, -53, -36, -62, -49, 2, 30, 17, 6, 5, 2, 67, 14, 14, 12, 47, 61, 27, 31, 28, -1, 25, 12, 53, 51, 40, 36, 12, 3, -16, -26, -67, -41, -16, 2, 13, -14, -21, -18, 39, 51, 41, 23, 12, 26, 11, 15, 28, 11, 42, 47, 30, 25, 22, 47, 24, 12, 3, -21, -38, -1, 2, 1, 0, 16, 19, 2, 28, 39, 49, 23, 20, 3, 49, 28, 35, 9, 27, 0, 18, 16, 45, 22, 38, 15, 2, 1, 19, 8, 8, -2, -12, 11, 7, -3, 47, 39, 13, 48, 13, 44, 59, 61, 38, 14, 10, -14, 11, 12, 56, 17, 6, 8, 28, 32, 45, 36, 38, 21, 8, 0, -12, 5, 3, 52, 47, 29, 8, 24, 44, 22, 14, 9, 12, -9, 37, 27, 25, 27, 0, -31, -39, -16, 45, 33, 22, 5, 8, 17, -12, -14, 29, 86, 40, 12, -23, -6, 18, -3, -13, 0, -42, -44, -22, 4, 14, 17, 41, 7, -7, 24, 43, 45, 42, -11, 13, 17, 2, 15, -19, 42, 85, 50, 15, 4, 59, 28, 38, 34, -17, -9, 20, 51, 24, 49, 38, 69, 47, 48, 68, 33, -19, 6),
  105 => (-1, -10, -2, -14, -14, -2, 12, 0, 11, -8, 12, -15, 5, -17, 19, -16, -3, 13, -6, 15, 29, 25, 11, 12, -6, 8, -14, 18, 11, 19, 11, -20, -17, -4, -17, -15, -4, 20, -19, -12, -4, 11, -17, -40, -42, -5, 35, 45, 6, 4, -9, -4, 2, -14, -13, 6, 20, 9, -16, -9, -18, 11, 9, 17, 17, -7, 11, 2, 3, 1, -28, -20, -41, -38, -8, -13, -17, -32, -56, 0, 41, 0, -1, -13, 10, -11, -20, -14, -5, -17, 2, -20, -6, -20, 0, 1, -25, -53, -35, -42, -47, -2, 38, 3, -51, -39, -37, 5, 58, 36, 19, 8, 19, 16, -20, 20, -4, -18, -1, 6, -34, 7, -43, -22, -32, -10, 22, 10, 12, 21, 13, -13, -36, -29, -2, 28, 3, 13, 16, 15, -2, 14, 1, 16, 0, -10, 8, -9, -33, 18, 29, 27, 3, 29, 15, 3, 14, 12, -11, -8, -31, -15, 0, 22, 6, 9, 11, -13, 9, 10, 3, -8, -5, 1, -28, -31, -2, 24, 23, 18, 31, 21, 6, 15, 22, 5, -31, -24, -18, -24, -9, 24, 27, 9, -10, -4, 10, 19, -18, -16, 1, -12, -35, -31, -51, -22, -30, -9, -5, 10, -17, -7, -10, 6, -13, -18, -8, -25, -41, -45, -1, 29, 28, 6, -18, -5, 8, -12, -1, -12, -13, -23, -89, -79, -70, -48, -39, -39, -31, -18, -28, -23, -44, -48, -14, 5, -16, -7, -33, 25, 15, 8, -19, -8, 10, -8, -14, -18, -45, -39, -79, -61, -46, -48, -75, -102, -28, -36, -32, -26, -54, -54, -10, 2, -22, -18, 5, 9, 29, 14, -1, 12, -6, -18, -2, 14, -2, -38, -71, -68, -34, -31, -89, -84, -16, -19, -15, -50, -72, -58, -18, 17, -13, -2, 11, 12, 24, 0, 6, 18, -11, 9, 16, 16, 26, -16, -56, -22, -42, -42, -40, -5, -3, -49, -4, -8, -55, -38, 31, 77, 50, 20, 26, -3, 24, 41, 4, -1, 13, -4, -9, 27, 85, 4, 10, -14, 16, -16, -1, 16, -2, 22, 4, 16, -9, -10, 23, 43, 10, 9, 1, 25, 19, 15, -17, 9, -18, -20, -4, 48, 122, 79, 74, 36, 66, 37, 59, 53, 48, 58, 25, 30, 17, 10, 54, 47, 32, 47, 12, 31, 25, -12, 13, 15, 13, -12, -56, 106, 113, 87, 58, 73, 55, 29, 39, 67, 65, 70, 37, 31, 7, 18, 8, 40, 51, 13, 17, 16, 39, 5, 3, 3, 3, 21, -7, 63, 41, 51, 37, 49, 53, 61, 19, 34, 7, 30, 11, -12, 5, 20, 7, 16, 50, 23, 10, -2, 31, 31, 19, -11, -2, -8, 1, 62, 12, 9, 24, 30, 46, -7, 15, 40, 35, 2, 10, -32, 11, 30, 9, 30, 12, 24, -5, 9, 45, 33, 11, 17, -15, 17, 16, 11, 33, 10, 32, 41, 53, 10, -10, 50, 66, 12, 1, 4, 3, 27, 11, 10, 5, 18, -18, 14, 29, 35, -20, 13, 20, 16, 9, 36, 41, 1, 5, 22, 62, 6, 34, 16, 14, -37, -50, -34, -33, 36, 6, -31, -11, -19, -12, 8, 7, 51, 2, 19, -11, -1, -6, 30, 7, -35, -25, -21, 31, -2, 8, -24, -11, -22, -43, 2, 2, 19, 12, -18, -17, -36, -41, -27, -64, 22, -9, 14, -17, 8, -32, -20, -58, -40, -82, -25, -23, 19, -4, -13, -21, -38, -39, -43, 6, 24, 24, -7, -6, -2, -43, -5, -36, -14, 9, -19, 18, -17, -5, -55, -44, -67, -50, -48, -39, -14, -26, -53, -30, -26, -52, -32, 3, 21, -3, -8, -15, -60, -14, 6, -25, 37, 10, 15, -17, -6, -24, -54, -14, -29, -20, 27, -15, -19, -55, -52, -18, 11, 5, -32, 18, 24, -4, -2, -5, -59, -42, -13, -25, 20, -19, 9, -19, 15, -17, -6, 10, -2, -22, -11, 1, -56, -41, -51, -40, -25, 24, 8, 35, 33, 19, 9, -39, -35, -23, -9, -12, 59, 15, 14, -10, -2, 0, 22, 9, -43, -36, -56, -45, -15, -49, -25, -32, 11, 3, 24, 12, 27, 45, -3, -39, -15, -19, 21, 0, 44, -6, -18, 2, 4, -3, 8, 49, -39, -5, -57, -28, -63, -63, -37, 10, -29, 9, 8, 49, 22, 32, 29, -6, -32, 10, 26, 42, 44, 8, 1, 9, -17, 28, 11, 10, -6, -12, -44, -32, -43, -53, -59, -32, -23, -36, -9, 8, 8, 44, 21, 2, -6, 3, 6, 17, 9, -12, 20, -2, -4, -20, 0, -18, 7, -29, -31, -48, -37, 5, -11, -12, -15, -24, -4, 12, -21, 1, 22, -11, -7, -19, 44, 14, 15),
  106 => (-4, 18, 5, -20, 19, -20, -4, -4, -11, -19, -14, 1, -20, 15, -5, 3, 17, 3, -26, -13, -32, -15, 12, 17, 14, -11, 5, -2, -14, -16, -6, 12, 13, -9, 7, 12, 1, -1, 21, -18, 8, 4, -15, -35, -31, -34, -55, -54, -50, -17, -47, 21, 17, 7, -14, -17, 5, -1, -13, 20, 13, -2, 12, 13, -10, 3, 15, -21, 6, -36, -55, -62, -89, -54, -27, -4, 5, 47, 20, 42, 35, -12, 21, -19, 2, -6, 1, 16, 12, -11, -15, 9, 14, -19, -16, 22, 23, -29, -31, -40, -58, -42, -52, -21, 4, -12, 23, 27, -57, 24, -7, -2, 12, -7, -10, -16, -20, 7, -1, -10, -5, -11, -14, 17, 15, -5, -4, -29, -31, -37, -47, 43, 34, 17, 40, 16, -53, -11, -7, 15, 17, 21, -10, 13, 4, 14, 15, -22, -16, -44, -44, -53, 25, -27, -20, -12, -60, -35, -49, 4, 19, 18, 35, 3, -29, -16, -14, -13, 6, -13, 5, -21, 13, -9, -18, -13, -25, -25, -36, -71, -10, 4, -24, -24, -30, -47, -31, 36, -3, 33, 39, -22, -1, 18, 17, 8, 19, 17, 1, 15, 18, -3, -29, -36, 9, -32, -70, -70, -13, -32, -26, -20, -22, -58, -26, -2, 17, 44, 50, 0, -16, -22, -19, -20, 5, 12, 18, -8, 4, 14, -33, 10, -5, -32, -36, -23, -7, -15, 14, -21, -42, -41, 20, 25, 37, 60, 11, -6, -15, -13, -13, 8, -14, -15, -10, -18, 8, 17, -13, -2, -27, -54, 9, -5, -9, -21, -37, -3, -44, -15, 19, 18, 2, 18, 7, -17, -6, -13, -46, -18, -15, 5, 13, -16, 7, 10, -31, -36, -33, -30, 10, 22, -32, -29, -34, -14, -28, 7, 34, 19, 15, 15, -6, -23, -26, -14, -10, 14, -8, 17, 4, -12, -4, -4, 17, -40, -53, -45, -18, -25, 16, 3, 14, -6, -3, 40, 22, 7, 61, 18, -5, -38, -52, -18, 5, -4, 16, 8, 2, -4, 15, 12, -17, -34, -51, -25, -20, -50, -49, -19, -45, -15, 33, 90, 5, 37, 48, 41, -28, 19, -35, -24, -23, -2, -6, 14, -16, 14, 12, -19, -52, -12, -29, -1, -8, -15, -47, -77, -28, 15, 61, 44, 8, 25, 23, -7, -26, -29, -53, -51, -23, 0, -13, -11, -5, 11, 2, -24, -25, -12, 22, 11, -24, 12, 7, -28, -19, 76, 89, 63, 11, 36, 5, -11, -29, -58, -56, -43, -22, 29, 2, -20, -2, -5, 28, 5, -11, -3, 23, 22, 38, 18, -8, -45, -25, 30, 77, 55, 43, 42, 26, -13, -33, -43, -49, -12, 31, 52, -2, -18, -19, -19, 17, 19, -23, 5, 43, 7, 46, -3, -34, -57, -37, 21, 31, 38, 3, 24, 16, -44, -87, -50, -84, -72, -45, 11, 9, 4, 19, 4, -14, -37, 13, -21, -15, -2, -1, -8, -64, -55, -15, 2, 46, 45, -3, 14, -24, -68, -83, -61, -52, -65, -22, 23, 6, -7, 20, -9, -31, -24, 20, 31, 9, 4, -13, -31, -23, -48, -2, 19, 50, 16, 19, -3, -34, -23, -16, -25, -43, -41, -39, 21, -2, -4, -12, 7, -13, 2, 23, 38, 36, 41, 21, -35, -13, -5, 22, 27, 47, 27, 1, -2, -18, -16, -17, -12, -47, -64, -69, -9, -1, 14, -3, 2, -12, -20, -14, -23, 10, -10, 20, -12, -42, -13, 18, 26, 19, 15, -9, -23, -8, -7, -15, -4, -43, -62, -33, -7, -14, 15, 10, -2, -5, 4, 3, -14, -48, -43, -44, -66, -42, -20, -3, 19, 1, 1, 20, -22, -32, -22, -41, -46, -93, -44, -27, -13, -17, -20, -11, 20, -6, -10, 20, -37, -39, -47, -27, -8, -9, 1, 19, 17, -17, -14, 20, 10, -33, -62, -80, -105, -91, -70, -19, 11, 19, -17, 11, -20, -18, 25, -7, -48, -41, -38, -50, 32, 17, 0, 6, 9, -7, -3, 21, 34, -28, -77, -108, -104, -89, -57, -20, -1, 18, -11, 17, 5, -27, -16, 18, -22, 5, 22, -35, 12, 4, 4, 1, 6, -10, 17, 11, 33, 26, -75, -70, -99, -49, -68, -20, 17, -4, 17, -14, 5, 10, -12, -10, -10, 5, 15, 23, 19, 13, -23, -6, 6, 0, -3, 28, 70, 14, -60, -56, -85, -70, -58, -20, -37, 2, 5, -18, 1, -19, -4, -14, 17, -31, 0, 10, 10, -3, 18, -14, 23, -7, -5, -14, 38, 73, -51, -64, -29, -58, -1, -3, 31, -10, -20, 11, 5, 4, 15, -21, -6, -42, 12, 2, 29, -8, 3, -20, -6, -22, 8, -15, 54, 58, -8, 4, -10, 22, 1, -11, -16),
  107 => (8, -19, 12, 13, 3, 18, -2, 14, 9, 6, -11, -20, 20, 1, -8, 30, 32, 27, -4, -29, -23, 7, -7, 6, 18, -14, 1, 18, -11, -8, 17, 8, -15, -19, -11, 0, -2, -8, -31, -1, 24, 32, 33, 1, 17, 32, 3, -13, -17, 27, -16, -20, 11, 10, 12, -7, -10, -15, -11, 17, 18, 1, -15, -2, 12, 4, 17, 26, -6, -10, 24, -12, -24, -25, 0, 9, 24, 33, 25, 42, 25, 12, -15, -4, -11, -3, 4, -14, -3, -3, 10, -21, -15, 14, -13, -25, -22, -19, -8, -11, 24, 17, 27, 19, 29, 36, 20, 34, 67, 19, 0, 13, -15, -19, -17, -14, -10, 6, 3, -47, 30, -4, -44, -24, -7, 0, -20, -16, 0, 24, 25, 23, 15, 21, 37, 35, 51, 26, -4, -8, 18, -2, -16, -2, 16, 9, 6, 1, 4, -33, -39, -37, 6, -7, -23, -1, -24, 26, 25, 19, 3, 40, 42, 10, -23, -31, -10, 15, -9, -10, 9, 16, -15, -1, 15, 5, 3, 4, -2, -32, 23, -4, -42, -12, -14, 25, 25, 12, -17, 33, 44, -9, -33, -13, 17, -15, 9, 15, 1, -15, 10, 17, 11, 6, -42, 25, 18, -17, 29, -4, -48, -18, 12, 26, 17, -7, -1, -6, 40, -10, -35, -4, -3, 12, 11, 5, 10, -3, 5, 3, -6, -13, -75, 24, -13, 4, 5, -3, -16, -13, 1, -7, 7, -25, 10, 26, 10, -16, -2, -17, 12, 20, 5, 9, -13, -16, -14, -11, -13, -28, -37, -9, 3, 4, 14, -16, -1, 31, 6, 3, -15, 0, 0, -8, 8, -6, 5, 24, -8, 18, 14, 1, 0, -16, -20, -20, -18, -18, 9, -14, 1, 10, -4, -33, 20, 5, 15, 1, 1, 1, 26, 30, 7, -17, -26, -19, 4, 8, -10, -7, -7, 17, -3, 9, 32, -46, -33, -8, -6, 21, -27, -31, 20, -2, -8, -4, -2, 10, 8, -5, -33, -57, -76, 0, -40, -8, -13, 18, 21, 19, -16, 58, 14, 13, 26, -3, -8, 11, -14, -19, -9, 12, -24, 9, -25, -6, 12, -14, -22, -33, -72, -50, -9, -31, -18, 2, 13, -3, 15, 18, 19, 7, 14, 5, 3, 12, 42, 26, -15, -41, 18, 38, -9, -6, -26, 0, -1, -25, -58, -64, -34, -11, -13, 12, -15, 0, 25, 3, 23, -16, 0, -12, -29, 16, 6, 15, -48, -27, -7, 5, 4, 1, -3, 2, -1, -9, -59, -27, -46, -15, -12, 19, 4, 8, 7, 50, 14, -21, -13, 4, 9, 49, 28, -9, -64, -45, 20, 28, -1, 12, 8, -13, -3, -31, -4, -40, -59, 10, -13, 3, 2, -7, 39, 33, -2, 11, 22, 28, 2, 40, 20, -6, -89, -35, 27, 1, 18, 10, -13, -24, 5, 8, -24, -28, -1, -17, 19, 0, 5, -7, 26, 29, 4, -2, 23, -2, 4, 47, 16, -64, -67, -16, 39, 18, 24, 28, -1, -13, -27, 8, -19, -69, 21, -6, 11, 20, -15, -14, 3, -26, -54, -40, -37, -1, 18, 52, -1, -49, -85, 19, 70, 19, 30, 30, -17, -52, -34, 9, -22, -51, 31, 23, 18, 13, -1, 18, -22, 6, -76, -45, 34, 0, 53, 52, -34, -100, -113, 30, 86, 22, 42, 31, -17, -62, -25, 14, -4, -17, -13, 31, 10, 4, -6, 5, -26, -3, -64, 10, 29, 15, 68, 29, -75, -113, -97, 21, 77, 36, 38, 50, 16, -45, -18, -40, -15, -14, -4, -9, -8, -18, 19, -10, 16, -10, -42, 30, 26, 25, 31, -29, -88, -137, -111, -7, 53, 31, 61, 56, 28, -46, -39, -59, -24, -26, -39, -8, 18, -6, -7, -18, 12, -11, 14, 84, 19, 14, 37, -49, -97, -125, -109, 5, 51, 31, 15, 68, 26, -12, -29, -43, -67, -69, -60, -33, 20, -7, -8, 20, 15, -13, 31, 35, 14, -1, 5, -53, -40, -88, -76, 1, 25, 2, 36, 9, 40, -31, -37, -45, -24, -59, -5, 4, 13, -20, -18, -12, -13, 6, 16, 39, -3, 4, -35, -100, -95, -108, -42, -12, -4, 7, 25, 22, 45, -27, -60, -54, -9, -57, -9, -20, 1, 10, -6, -1, 16, 9, 19, 20, -1, -34, -67, -121, -138, -128, -60, 28, 27, 48, 57, 18, 32, -43, -85, -66, -46, -40, -6, -38, -3, -12, 3, 15, -8, 21, 15, 3, 7, -36, -47, -90, -113, -106, -63, 11, 24, 15, 10, 32, 17, -47, -50, -39, -12, -5, 7, -31, 18, 3, 20, 11, -11, 13, 13, -9, -14, -23, -20, -57, -63, -79, -42, 5, 46, 45, 1, 27, 58, -16, -25, -36, -39, -22, 20, -14),
  108 => (16, -13, 7, 20, -8, 17, -14, 18, -19, -12, -18, -8, 0, -10, 19, -25, -8, -4, 17, 5, 6, 8, -5, 19, -20, -19, -2, 9, 15, 16, -10, 3, 13, -6, 8, 12, -16, 0, -15, 5, 27, 21, 28, -20, -7, -5, -5, 14, 25, 25, 4, 49, 13, 16, -19, 3, 3, -5, -11, 0, 7, -19, 7, 3, 2, -40, 7, -21, 6, -1, -14, -28, -49, -36, -47, 23, 1, 16, 28, 28, 42, 11, -6, -17, 3, -20, -16, 8, -1, -11, 8, -10, -37, 12, -15, -37, 3, -26, -47, -44, -23, -48, -8, -22, -7, -15, 3, 15, 44, 27, -11, 1, 10, 12, -14, 2, 13, -9, -2, -38, 7, -13, -24, 7, 5, -1, -16, 3, -41, -52, -65, -28, -26, -5, 8, 24, 25, 13, -6, -6, 2, 20, 6, 1, 12, 11, 10, 3, -25, -71, -50, -26, -51, -25, -46, -28, -10, -20, -51, -46, -28, -11, 39, 49, -10, 31, -13, -13, -8, -20, 12, -15, 2, 2, 5, 4, -28, -24, 20, 16, -10, -4, -33, 12, -17, 9, -8, 0, -13, 14, 54, 8, 35, 19, 7, 17, 15, 10, -10, 12, 16, 1, 8, 2, -49, 39, 55, 34, 13, -1, -4, 12, 33, 28, 15, -17, -26, 10, 7, 28, 16, 0, -3, 2, 14, 6, 11, -1, 9, -15, -26, -45, -22, 13, 22, 13, -6, 23, 0, -5, 5, -5, 9, 1, 7, 6, 37, 34, 38, 11, 8, 11, 11, -10, -16, -20, 18, 4, -10, -49, -57, -1, 11, 18, 21, 18, 6, -6, 52, 11, 12, 20, -22, -8, 12, 10, 10, -7, -36, 3, 10, 14, -19, -10, -11, -24, -73, -47, -10, -35, -29, -4, 6, -16, -2, 4, 10, 6, -13, 18, -7, 4, -5, 25, 0, 5, -31, -43, -5, -2, 3, -6, -16, -10, -46, -62, -65, -70, -72, -50, -7, -2, -42, -6, -7, -11, -7, 10, 4, -5, 20, 14, 5, -11, -46, -26, 6, 1, -6, 19, 16, 45, -20, -35, -66, -101, -61, -30, -1, -26, -31, -12, -27, -16, 2, -10, 13, 9, 0, 13, -21, -41, -57, -42, -12, -1, -12, -7, 6, 50, 13, -27, -29, -60, 0, 17, 0, 4, 19, -14, -7, -36, -14, 15, 11, 13, 19, 3, -17, -27, -34, -11, -4, 7, -2, -16, 14, 28, 31, 33, 1, 31, 27, 37, 39, 29, 20, 13, 17, -21, -30, -10, 14, 45, 17, -41, -34, -2, -2, 14, 0, 9, -16, 2, 1, 13, 44, 43, 33, 26, 8, 50, 50, 21, -12, 16, -40, -52, 7, 46, 38, 23, 10, -11, -24, -42, -11, 24, 20, -4, 11, 18, 1, -10, 33, 14, 18, -15, -6, 28, 75, 36, -15, -10, -34, -45, -24, 11, 19, 18, 1, -30, -24, -25, -3, 30, 17, -16, -6, -15, -30, 21, 20, 18, 8, 12, 20, 65, 80, 25, -16, -21, -56, -18, 1, -2, 10, 41, -18, -9, -3, -7, -1, 37, -16, 15, -11, -4, 2, 29, 28, -4, -16, 7, 36, 71, 33, 18, -11, -29, -68, -71, -1, 9, 38, 55, -1, -4, -6, -9, -4, 21, -7, -11, 2, 1, 32, 28, -20, -11, -69, -49, 16, 20, 29, 5, -20, -63, -125, -97, 3, 13, 24, 35, -4, -26, -3, -22, -16, 27, -2, 3, 18, 12, 50, 11, -5, -41, -84, -52, 19, 35, 26, 29, 3, -75, -84, -113, 10, 24, 22, 41, 23, -33, -42, -46, -43, 6, -19, -8, 7, -2, 30, -7, -48, -51, -51, -35, 32, 64, 23, 35, 29, -52, -85, -93, -55, 16, 13, 33, 12, 7, -23, -16, -19, 27, -15, 8, 17, 4, -9, -22, -71, -85, -86, -63, -25, 15, 9, 65, 25, -74, -91, -83, -14, 51, 17, 10, 11, 52, 14, -4, 11, 72, -15, -1, 0, -5, -9, -37, -45, -77, -103, -73, 2, 42, 10, 21, 21, -42, -82, -73, -38, 2, 22, -16, 32, 37, 12, 6, 29, 72, 12, -7, 9, 13, -15, -9, -53, -36, -56, -24, 20, 43, 37, -31, -23, -49, -71, -42, -50, -23, 22, -3, 26, 21, -7, -19, 33, 48, -5, 13, 16, -6, -15, -23, -27, -54, -32, -45, 34, 42, -19, 8, -49, -28, 3, -1, -30, -16, 16, 15, 24, 7, 3, -24, -22, 26, -5, -13, -6, -8, -8, 13, -13, 14, -29, -34, 2, 36, 21, -7, 0, -22, 14, 12, -1, 4, -8, 12, 11, -26, -22, 23, 17, 1, -3, 5, -17, -13, 19, 16, 6, -2, -23, -9, 20, -6, -7, 20, 14, -4, 8, 39, 30, 49, 17, 6, 31, 14, -15, -31, 3, 18),
  109 => (-12, -15, 0, 17, -10, 7, 10, -15, 15, -16, 19, -17, 17, -12, -20, -23, -3, 15, 21, 5, -44, -33, 3, -1, -15, 6, -16, 12, -9, -1, -8, 0, 5, -7, 14, 0, 19, 9, -13, 16, -39, -16, -15, -4, -7, 11, 11, 26, -30, -20, 2, -13, -12, 20, 14, 20, -6, 15, -12, 12, -7, 7, 0, 18, 1, -4, -2, -26, 20, 23, 7, 2, 1, 21, -12, -27, -11, 3, 20, 20, -2, 5, -6, 17, 6, -9, -7, -20, 6, -14, -1, 12, 26, 4, 10, 13, -6, 8, -15, 12, 19, 17, 18, -12, 6, -17, -2, -9, -25, -30, 2, -19, 14, 7, 14, 5, -20, 18, -8, -2, 14, 43, 37, -23, -22, -11, -8, -3, 11, 27, 25, -8, 1, 16, 0, -18, 2, -32, 15, 4, 5, 10, 4, -13, -1, -8, -11, -1, 14, 52, 7, 13, -47, -25, -60, -17, 29, 10, 9, -9, 11, -11, 4, -39, 28, 20, 19, 5, -5, 7, -12, -6, -6, 7, 1, 12, 70, 27, -7, -27, 10, 0, -17, 17, -18, -17, -4, -1, -1, -10, 7, -13, -11, 38, 2, -19, -11, -10, 12, -16, -14, -13, -23, 37, 6, 13, 8, 38, 26, 35, -16, 12, 4, -12, -41, -19, -21, -13, -9, -4, 5, 48, 15, 16, -16, 9, 12, -18, -3, -6, -25, 40, -22, -19, 24, 49, 34, 21, -26, -10, -9, -12, -14, 10, 13, 13, 1, 7, 2, 36, 17, 17, 7, 8, -1, -19, -19, 12, 19, -19, -29, -6, 14, 17, 8, 6, -11, 0, 10, -16, -14, -1, 7, -15, -23, -1, 32, 48, 15, -36, -11, 17, -3, -19, -17, 0, 28, -2, 8, -14, 24, 3, -32, 6, 16, -12, -19, -16, -39, -29, -26, -3, -39, -4, -3, 44, 41, -28, 17, 0, 16, -13, -16, 31, 6, -15, 15, 17, -4, 18, -24, 11, 17, -14, -18, -25, -22, -28, -30, -3, -27, -12, 17, 26, 16, 11, -6, -5, 19, 18, 8, 47, -24, 11, 25, -6, -10, 16, -33, -20, -4, -31, -39, -22, -15, -29, -26, 8, 12, 3, 42, 44, 31, 8, -2, -9, 7, 14, 33, 70, 36, 25, 8, 4, -27, -28, -43, -34, -20, -30, -50, -56, -18, -32, -30, -17, 26, 21, 27, 32, 46, -15, -19, 20, 17, 14, 24, 34, 8, -21, -48, -62, -24, -41, -56, -77, -29, -59, -52, -12, -38, 3, -9, 23, 43, 42, 26, 35, 22, 12, -8, 19, -14, 7, 35, 11, -21, -45, -87, -85, -81, -89, -107, -101, -48, -31, -28, -2, 31, 28, 52, 40, 7, 24, 15, 56, 32, 6, 14, -18, 4, -14, -18, -34, -31, -97, -100, -104, -93, -96, -75, -56, -5, 4, 8, 41, 65, 54, 28, 12, 19, 2, 16, 5, 17, 47, -4, -2, -17, -10, -31, -5, -31, -71, -37, -57, -22, -6, 13, 48, 64, 78, 67, 58, 48, 47, -2, -16, 16, -18, 13, -17, 14, 14, -15, -10, -1, 19, 5, 17, -6, 25, 3, 16, 42, 66, 67, 50, 36, 49, 42, 42, 35, 11, 16, -11, 34, -13, -19, 16, -9, 37, 9, -10, 16, 13, 28, 32, 63, 36, 22, 22, 58, 41, 40, 27, 15, 25, 48, 13, -1, -13, 22, 21, -10, -25, -12, 13, 22, -27, -7, 2, 19, 2, 30, 41, 57, 34, 51, 37, 39, 49, 63, 40, 23, 13, 15, -17, -30, 5, -15, -48, -40, -44, 1, 4, -15, 5, -4, 12, -10, 2, 9, 34, 52, 71, 42, 43, 37, 35, 82, 45, 28, -21, -15, -36, -14, -26, -41, -25, 0, 3, 20, -14, -15, -1, -7, 6, 5, 11, 27, 16, 2, 41, 26, 38, 5, -7, -13, -17, -3, -46, -17, -29, -10, -18, -57, -6, -11, -14, 7, -1, -2, -26, -17, -1, -7, 10, 60, 23, 47, 36, 24, 37, -14, 4, -23, -38, -26, -7, -16, -19, -6, -46, -29, -54, -27, -3, -19, -34, -15, 0, 6, -2, 11, 18, 34, 12, 12, 13, -11, -42, -49, -69, -62, -48, -72, -45, -45, -29, 25, -34, -37, -32, -13, -18, -54, -19, -18, 0, -17, -11, 8, -6, 6, 17, 50, -1, -13, -7, -31, -84, -76, -68, -44, -45, -52, -52, 11, -14, -24, -49, -27, -32, -49, -37, 12, -5, 19, -9, -16, 2, 2, -34, -2, -2, -13, -33, -59, -57, -54, -42, -75, -36, -68, -29, -37, 1, -50, -17, 0, -25, -30, -15, 1, 2, 10, -2, -3, -5, -1, -30, -19, -14, 3, -43, -22, -49, -21, -42, -47, -44, -44, 1, -9, -49, -10, 12, -21, -23, 6, -15, -2, 3),
  110 => (-4, 3, 14, 12, -16, -10, -2, -19, 11, -10, 11, 6, 16, -8, 23, -22, 15, -8, 17, 14, 44, 24, 10, 4, -17, 8, 17, -17, -13, 4, -12, 0, -14, 18, 15, 7, 4, 17, -7, -3, -6, 23, 28, 3, 4, -9, -13, -1, 2, 12, -7, 27, 15, 3, 9, -12, -9, 19, 17, 5, -14, -4, 5, 7, -8, -1, 12, 0, 45, 45, -1, -10, -22, -63, -41, -38, 16, 17, 52, 50, 19, -6, -8, 4, -21, -2, -13, 1, 15, 12, 12, 8, 13, -11, 24, 49, 55, -18, -40, -36, -71, -60, -23, -29, -22, 49, 11, 31, 45, 35, 11, 16, 17, 20, 12, 16, 13, 0, -1, 14, -16, 32, 39, -5, -33, -26, -37, -41, -62, -48, -12, -5, 15, 29, 28, 38, 44, 25, 1, -6, 3, -5, -1, 8, 17, -8, 28, -4, -11, 12, -5, -79, -40, -13, 21, -15, -36, -30, -18, -17, 30, 28, 21, 20, 30, -16, 1, -20, 8, -6, 19, -6, -14, -2, 31, -34, 43, 16, -64, -75, -13, -1, 24, -12, -36, -33, -17, 4, 12, 39, 39, 30, 29, -3, 3, -14, -8, -20, -14, -6, -14, 13, 42, 26, 63, -18, -107, -73, -18, 0, 6, -7, -40, -45, 7, 16, 18, 24, 16, 28, 17, 2, -12, 15, 9, 14, 6, 2, 6, -16, 22, 54, 0, -35, -35, -54, -14, 7, -6, -39, -27, -41, 11, 31, 45, 35, 33, 34, 46, 19, -36, -9, -12, -8, -3, -18, 13, -1, 63, 50, 29, 18, 30, -26, -15, -18, -11, 2, -28, -30, 12, 23, 30, 9, -13, -14, 58, -6, -17, -7, -17, 14, -14, 5, -13, -11, 80, 34, 7, 40, 17, -16, 14, 32, -7, -10, -27, -29, 10, 20, 24, 14, -14, -20, 13, 1, -1, -21, 0, -9, -13, 2, 12, -13, 39, 2, 23, 47, -23, -14, 1, 4, -27, -25, -30, 17, 31, 25, 41, 31, 27, 13, 9, 4, 10, 0, -14, 11, -14, -15, -48, -3, -12, 26, 47, 24, 1, -29, -3, -29, -27, -2, -7, 28, 70, 7, 33, 8, 18, -14, -34, -16, 37, 52, -12, 2, 6, -4, -30, -25, -5, 22, 35, 38, 13, 28, 2, -5, 13, -9, -16, 70, 48, 19, 31, 21, 16, -15, -3, -30, -21, 46, 13, -8, 2, -1, -39, -6, 20, 42, 32, -3, 0, 29, 22, 10, -5, -34, -17, 60, 31, 7, 6, 10, 33, -26, -29, -4, -3, 43, -9, -7, -6, 1, -20, 16, 40, 47, 33, 36, 4, 0, 35, 16, -9, -16, 7, 77, 29, 29, 7, 19, 27, -28, -19, -22, -25, 57, -18, 12, 8, 5, -27, 18, 35, -7, 35, 20, -7, 9, 17, 22, -18, -19, 6, 52, 28, 18, 14, -13, -6, -44, -37, -45, -5, 54, 10, -9, 7, 15, -62, 7, 3, -28, 16, 0, -12, -12, 18, -2, -25, -69, 20, 54, 26, 20, 4, 20, -16, -24, -42, -48, 9, 58, 12, -16, -12, -16, -40, 1, -11, -16, 8, -19, -58, 6, 34, 12, -38, -70, -32, 18, 35, 36, 28, 9, 37, 35, -26, -54, -10, 50, 10, 14, -10, 2, 9, 18, -5, -26, -7, -52, -62, 6, 9, -43, -67, -97, -46, 43, 39, 22, 10, 5, 15, 6, -12, -57, -52, 51, -15, 15, -13, 9, 6, 24, -12, -17, 23, -38, -34, 21, 2, -66, -109, -114, -57, -11, 24, 7, -6, 27, 20, 21, -41, -76, -77, 36, 6, -15, 11, -11, -16, 64, 24, 36, 33, -28, -8, -11, 15, -44, -116, -103, -54, 2, 6, 7, 16, -4, 16, -16, -21, -97, -70, 16, -12, 7, -6, 18, -5, 63, 26, 25, 5, 5, 1, 26, -14, -48, -75, -38, -13, 22, 37, 67, 46, 49, 63, 28, -27, -120, -63, 21, 15, 20, -16, -17, 13, 61, 72, 55, 16, -65, -50, -10, -10, -35, -61, -12, -4, 4, 13, 20, 53, 58, 69, 32, -44, -143, -94, -30, 3, -2, 3, -11, -14, 26, 27, 31, -5, -41, -36, -12, -33, -64, -45, -19, 0, 26, 31, 12, 27, 28, 4, -3, -35, -106, -86, -51, -2, -12, 1, -11, -13, 27, 24, 36, 18, 12, -14, 10, -1, -62, -94, -65, -23, 26, 8, -6, 24, 10, -3, 6, -33, -65, -33, -1, 12, 2, -13, -16, -1, 21, 32, -2, -5, 2, -25, -25, -5, -33, -96, -64, 11, -10, 7, 13, 36, 35, -3, 4, -82, -44, -40, 18, -10, 0, 11, -18, 0, 24, 19, -36, -36, -20, -5, 7, 9, -18, -56, -29, -26, -26, -24, 38, 30, 3, 17, -19, -59, -80, -29, -6),
  111 => (18, -5, 10, -20, -12, 7, -10, -10, 11, -4, -7, 5, -6, 0, 10, 2, -2, 16, 7, 4, -24, -21, -8, 2, 8, 10, 0, -10, -12, 1, 1, -3, -10, 3, -1, 3, 20, -12, -7, 4, -26, -5, -24, 0, -8, -12, -12, -20, -11, 6, -41, 32, 16, -15, -4, -12, 4, -3, -5, -5, -18, 0, 2, 5, -18, -17, 0, -30, -3, -14, -39, -13, -35, -27, -31, -18, -39, -31, 13, 2, 22, 26, 10, 0, -4, 6, -11, 5, 0, 11, -18, 1, 2, -30, -42, -46, -76, -48, -53, -28, -29, -37, -7, -38, -13, -36, 7, 4, 5, -32, -15, 16, -1, 19, -4, 1, 15, -14, -9, 16, -25, -78, -78, -16, -6, -3, -19, -16, -40, -28, -22, -36, -33, -34, 6, -7, -22, -41, -5, 10, -10, 17, -2, -4, 20, 19, 11, -27, 3, -2, -20, -34, 14, -19, -46, -26, -33, -25, -37, -31, -17, -30, -27, 3, 2, -29, -12, -17, 17, -4, 8, 8, -10, 3, -23, 6, 28, 10, -31, -23, 19, -30, -35, -10, -43, -28, -38, -47, -4, -29, -36, 26, 28, 23, 15, -3, 20, -6, 17, -18, 19, 16, 1, 18, -10, -57, -22, -4, -11, -20, -13, -9, -15, 1, -19, 5, -2, -9, 12, 6, 10, 34, 17, 20, 11, 19, 15, -13, 0, 18, 14, -1, 7, 9, 17, 16, 18, 0, 7, -7, 8, 7, 3, 27, 25, 25, 50, 45, 28, 52, 39, 61, -7, 10, 12, -14, -4, 1, -5, 44, 50, 22, 59, 53, 49, 42, 15, 4, 9, 22, 28, 24, -3, -5, 41, 36, 51, 37, 29, 42, 4, -11, 9, 1, 11, 47, 27, 83, 63, 57, 29, 27, 53, 51, 7, -3, 2, 16, 31, 19, 35, 32, 36, 3, 28, 7, 24, 50, -7, -14, 6, 1, -19, 65, 72, 99, 60, 57, 34, 28, 21, 29, 33, 1, 23, 17, 7, -10, -16, 5, 33, -25, -7, -11, -2, 8, 7, 3, 0, -12, 8, 64, 35, 9, 40, 44, 39, 52, 31, 24, -8, -8, 2, -20, -12, -11, -38, 9, 1, -21, -5, 1, -32, 12, -19, -19, 3, -17, -34, 61, -20, 8, -3, 9, -5, -14, -81, -42, -72, -61, -55, -38, -8, -28, -20, -7, 1, -9, 35, 17, 0, -8, 20, 17, 0, -19, 4, 21, -9, -66, -57, -48, -80, -102, -96, -44, -31, -48, -47, -15, -35, -27, -10, -22, -17, 1, -11, 2, -23, -10, 9, -13, -16, 11, -19, -42, -40, -35, -67, -70, -65, -61, -74, -17, -14, -28, 4, -21, -22, -20, -1, -11, -6, -22, 9, 14, -28, -10, 18, -16, 0, 0, -13, -50, -75, -79, -102, -90, -19, -38, -32, -14, -8, -25, -27, -32, -30, -14, -7, -13, -9, -6, -15, -18, -18, 8, -9, -8, 17, -10, -30, -44, -62, -65, -75, -59, -36, -19, -69, -30, -55, -49, -49, -55, -46, -44, -4, -18, 10, -28, -28, -12, -17, -25, -19, 10, 2, -9, -18, -40, -71, -61, -51, -58, -78, -73, -79, -70, -18, -6, -19, -16, -26, -8, -17, 15, -15, -9, 4, -10, -25, 38, -10, -11, 1, 7, -57, -51, -48, -44, -85, -78, -39, -15, -65, -21, -2, 21, 14, 4, -5, -19, 37, 8, -1, -20, 0, -20, -6, 42, -6, 5, -5, 19, -11, -57, -45, 19, -8, 4, 15, 30, -34, -18, 0, 1, 11, 20, 20, 30, 33, 17, -7, 21, 22, -11, 7, 32, -9, -14, -17, -16, 12, 13, -38, 42, 40, 18, 31, 13, 0, -30, -2, -9, 38, 43, 18, 19, 25, 18, 17, 17, 28, 7, 4, 33, 4, -11, -10, -13, 18, 12, -21, 14, 36, 21, 6, 8, 4, 26, 61, 38, 61, 27, 29, 9, 28, 27, 30, 14, -43, -46, -26, 44, 8, 16, 10, -20, 13, -2, 4, 27, 14, 1, -13, -6, 29, 54, 41, 46, 49, 24, 2, 48, 42, 41, 18, -33, -75, -45, -36, -1, 4, 15, 10, 13, -1, 10, 45, 2, 0, 5, 0, -13, 4, 12, -1, 4, 18, 25, 18, 5, 0, 37, 20, -7, -46, -37, -27, 34, 7, 11, 6, -3, 14, 0, 10, 8, -15, -2, 19, 2, 16, 56, 21, 7, 3, -10, 6, -45, -63, -28, -14, 9, -11, 3, 36, 48, -3, -10, -9, 5, -10, -36, -1, 44, 30, -1, 4, 38, -8, 18, 16, 15, 2, -11, -21, -34, -56, -70, -37, -10, 9, 17, 40, 40, -19, -6, -2, 0, 15, -10, -2, -23, -10, 8, -3, 24, -19, -40, -53, -43, -50, -30, -37, -34, -10, -28, -1, -38, -14, 25, 31, 69),
  112 => (-19, 1, 16, -2, 10, 7, -12, 10, -19, 15, -6, -12, -18, -19, 0, 1, 4, 24, 1, 8, 9, -25, -30, 6, 12, -6, 11, -18, -13, -3, 2, -20, -21, 0, -3, 16, -17, -14, 13, -38, 9, -3, -2, 42, 36, -11, -9, 9, 43, 37, 4, -18, -11, 1, 9, 12, -10, 15, 2, 16, -7, -5, 5, 4, 3, 25, -9, 5, -12, -5, 9, 33, 48, 20, 3, 15, 10, -12, -32, -15, 18, -22, -12, -12, -12, -6, 4, 10, -15, -7, -20, 5, 0, -21, 40, -19, -2, -42, -15, 22, 33, 33, 0, -4, -12, -38, -41, -40, -37, 6, 18, -20, -16, 7, -18, -13, 15, -11, 20, 1, -12, 3, -21, -32, -10, -38, -15, 24, 26, -15, -24, -45, 0, -3, -17, 4, -7, 5, -5, -3, -5, 8, 20, 13, 14, 14, -12, 6, 19, -29, -41, -41, -74, -71, -6, 18, 36, 6, -32, -19, -20, -26, -9, -11, -61, 19, 19, -2, 8, 20, -20, 7, 11, -19, 10, 1, -8, -6, -46, -67, -43, -35, -6, 7, -10, -23, -37, -35, -38, -35, 16, 4, -36, 6, -6, -4, 5, 9, -3, 12, 9, 7, 6, -21, 10, -14, -63, -69, -41, -27, -8, -26, -4, -22, -60, -37, -2, -7, -27, 3, -18, 10, -8, 3, 17, 10, 12, 13, 2, 6, -35, -13, -30, -55, -32, -52, -43, -18, -32, -38, -33, -23, -37, -30, 30, -10, -45, -37, -11, 1, 1, 16, 5, -5, -1, -11, 19, -15, -16, -54, -45, -42, -46, -20, -46, -24, -68, -48, -56, -15, 0, 5, 1, -55, -60, -29, -20, -37, 45, 10, -16, 14, -1, -13, -18, -11, 16, -55, -63, -70, -62, -57, -61, -50, -53, -4, 8, 5, -6, -2, -9, 5, 11, 26, 12, -27, 57, -4, -11, -5, -18, 13, -12, 26, 9, -54, -65, -48, -65, -26, -12, 9, -7, 19, 38, 30, -10, -22, 22, -2, 33, 35, 37, 12, 23, 19, 1, -19, -9, -7, -18, 9, -18, -41, -20, -28, -38, -4, 5, 4, -1, 24, 10, 43, 23, 30, 41, 24, 33, 47, 53, 12, 16, 3, 17, 9, -5, 8, -5, 36, -36, -26, -13, -6, -11, 1, 28, 32, 36, 30, 50, 49, 50, 45, 31, 43, 21, 47, 31, 26, 50, -14, -15, -8, 20, -14, 11, 47, 22, 19, 10, 2, 30, 55, 35, 42, 47, 32, 54, 32, 12, 23, 23, 19, 39, 38, 51, 38, 18, 46, -7, 12, 11, -4, 16, 60, 41, 33, 45, 47, 22, 48, 32, 7, 38, 44, 42, 40, 20, 4, 31, 1, 7, 23, 13, 11, 22, -19, -17, -2, 18, -9, 34, 58, 28, 26, 37, 20, 43, 36, 24, 54, 18, 29, 41, 5, 28, -12, 2, -8, 23, 36, -5, -1, 4, -13, 2, -11, 13, 3, 10, 43, 38, 59, 44, 44, 46, 48, -12, 26, -15, 4, 1, 29, 23, 18, 11, -19, 27, 11, 25, 9, -44, 33, -13, 15, -18, 15, 35, 23, 20, 25, 42, 4, 44, 16, 1, 19, 19, -23, 25, 10, -9, 2, -16, -7, -22, -22, -22, -32, -68, 15, -19, -14, 3, 12, 13, 29, 19, 35, 45, 38, 19, 62, 19, 24, -20, -11, 5, -1, -10, -8, -8, -13, -2, -28, -41, -8, -26, 34, 12, 20, 4, 5, -1, 19, 14, 10, 23, 28, 50, 26, 28, 11, -29, -44, -7, -25, -3, 3, -36, -9, -33, 0, -24, -2, -24, 29, -4, -2, -13, -20, 19, 19, 12, -7, -64, -26, -27, -25, -24, 14, -39, -22, -23, -25, -31, -20, -25, -16, -51, -35, -24, -8, -14, -24, 13, 3, -8, -13, 25, 3, -3, -29, -61, -23, -18, -36, -41, -47, -59, -72, -70, -78, -70, -67, -16, -54, -62, -65, -69, -44, -49, 10, -20, -16, 9, -17, 28, 27, -29, -46, -55, -51, -47, -60, -23, -76, -41, -50, -44, -26, -33, -42, -39, -51, -38, -80, -81, -14, 8, -9, -12, -5, -10, 20, 11, 11, -56, -36, -28, -26, -62, -74, -27, -76, -59, -44, -54, -39, -31, -31, -50, -11, -22, -40, -44, 16, -2, 11, 12, -15, -15, 20, -14, 4, -6, -51, -62, -50, -72, -48, -42, -66, -41, -28, -41, -17, -29, -51, -61, -14, -23, 17, -41, -13, -4, -6, 18, 5, 1, -18, -13, -11, -35, -24, -58, -29, -44, -47, -36, -16, -3, -41, -34, -20, -33, -28, -7, -42, 6, -19, -1, -45, -16, -16, 0, -4, 14, 5, 2, 0, -8, 1, -48, -47, -31, -73, -34, -33, -50, -35, -46, -62, -51, -64, -40, -57, -25, -47, -3, -35, 17, 16),
  113 => (-4, 20, -1, 18, 7, -16, 19, 18, 18, 3, -9, -5, -7, -12, 1, -32, 0, -10, -29, -13, -1, -11, 16, -1, 4, 8, 17, 15, -21, -20, -1, 14, 19, 5, -16, -9, 19, 3, 7, -1, 23, 8, 17, -35, -10, -9, 28, 18, 16, 37, 34, 15, -11, 10, 15, 18, -3, 21, -16, -8, 19, -15, -5, -3, 1, 19, 0, -32, -19, -13, -11, 12, -13, -13, 20, 1, 54, 75, 62, 3, 0, 14, 0, -13, -20, -11, -2, -1, 7, -8, 3, -5, -7, -4, -9, -17, 0, 5, 17, -7, -36, 2, 7, 43, 18, 8, 31, 27, 0, -9, -14, 2, -6, 19, 10, 11, -4, 11, -13, 21, 7, -22, -4, -9, -11, -20, -16, -11, -15, -15, -2, -17, 14, 6, 2, 3, -1, 7, -19, -9, 9, -4, -11, 0, 4, 21, -5, 10, -28, -35, -4, -4, -16, 3, -8, -7, -39, 17, -8, 20, 23, 50, 7, -15, -3, -2, 16, -19, 15, 5, -15, 9, -9, 6, 5, 3, -24, -20, -28, -28, -17, 15, 26, -7, -7, 15, 7, 24, 30, 35, -1, -21, 3, 47, -15, -9, -16, -17, 8, 10, 14, 4, 20, -24, -2, -13, -40, -46, -18, -17, 10, 10, 15, -11, 7, -6, -3, -6, 1, -18, -12, 12, -16, 11, -18, 4, -2, -13, 2, -3, 30, -40, 9, -32, -29, 0, -37, -28, 9, 13, -19, -11, -31, -19, -36, -46, -54, -63, 18, 30, 19, 12, -18, 1, -14, 11, 9, 5, 18, -14, -21, -19, -42, -20, -31, -42, -15, 24, -2, -46, -66, -22, -36, -22, -71, -52, -17, 24, 28, 7, 18, 14, -10, -20, 1, -25, -27, -38, -28, -35, -30, -17, -27, -24, -29, -2, -13, -47, -52, -29, -39, -44, -76, -60, -23, 5, 11, 2, -1, 15, -10, -6, -20, -13, -38, 23, -43, -18, -23, -42, -62, -60, -22, -74, -32, -46, -45, -62, -65, -72, -89, -58, -9, 28, 4, 28, 13, 0, -16, -2, -5, -23, -26, 4, -21, -33, -11, -19, -11, -37, -60, -66, -35, -26, -36, -30, -47, -18, -52, -64, -4, -24, 38, -2, 14, 20, -13, -17, 4, 7, -10, 6, -49, -25, -34, -3, -42, -31, -23, -42, -1, -1, -21, -19, -20, -6, 13, -18, -7, 22, 11, -10, -2, 7, 19, 18, -14, 14, -8, -14, -41, -81, -18, -13, -27, -46, -23, -46, -8, 37, -25, -60, -31, 12, 4, 5, 52, 46, 32, 21, -1, 15, -19, -15, 0, 16, 13, -22, -25, -20, -43, -43, -24, -23, -32, -38, 8, -6, -18, -10, 15, 27, 8, 27, 22, 65, 54, 50, -20, -8, 1, 20, 7, 23, 33, -2, 4, -17, -8, -3, 6, -11, 2, -44, -8, 15, 22, 26, 31, 5, 34, 59, 72, 40, 34, 30, -7, 18, -9, 15, 27, -3, 45, 55, 9, 0, -4, 53, 54, 18, -3, -4, 55, 38, 40, 13, 28, 31, 42, 63, 39, 40, 58, -5, -19, 2, -10, 10, 17, -4, 44, 26, 39, 19, 57, 65, 58, 66, 17, 18, 48, 57, 23, 30, 25, 44, 49, 35, 38, 59, 51, 51, 10, 14, -3, -15, 43, -5, 40, 59, 28, 36, 73, 103, 83, 61, 20, -20, 26, 39, 52, 5, 20, 16, 16, 45, 29, 20, 34, 52, -7, -8, -9, 4, -17, -11, 25, 63, 19, 22, 36, 24, 63, 95, 74, 10, 26, 20, 24, 47, 24, -16, 44, 58, 25, 1, 9, 56, 19, 1, 5, -3, 8, 34, 21, 46, 26, 50, 37, 31, 33, 49, 54, 40, 44, 16, 6, 15, 1, 1, 54, 50, 18, 33, 33, 33, -12, 11, 11, 0, 19, -4, -2, 51, 32, 18, 49, 10, 39, -4, 48, 49, 28, 54, 10, 28, 19, 22, 67, 11, 5, 7, 32, 74, 12, -7, 16, 4, 10, 15, -5, 28, 39, 34, 46, 22, 3, 45, 28, 49, 52, 26, 29, 43, 43, 61, 0, -18, -32, 14, 63, 86, -8, -14, 7, -3, -5, 22, 18, 30, 63, 27, 31, -5, 37, 26, 39, 27, -9, -17, 22, 31, 31, 29, 26, 24, 8, 7, 51, 79, -18, -11, -9, 0, 43, 29, 38, 1, 25, 15, -8, 8, 4, -10, 15, 41, 10, 9, 21, 20, 15, 23, 30, 11, 12, 35, 48, 73, -16, -16, -9, 3, 11, 44, 64, 17, -2, -33, -44, -59, -48, -56, -44, 2, 13, -11, 14, 24, 27, 24, 26, -1, 48, 44, 69, 83, 19, -2, -15, 16, 4, 22, 1, 57, 50, -5, 0, -34, -42, -17, -6, 27, 29, 18, 44, 78, 25, 44, 41, 36, 25, 58, 58, 20),
  114 => (-6, 6, -4, 5, -13, -2, -17, -18, 16, -13, 14, -10, -4, -2, 0, 8, 74, 57, -4, -34, -8, -20, 1, 2, -18, 12, -16, 6, 5, 14, -20, 9, -7, -14, 0, 20, 20, -20, -3, 51, 34, 41, 17, 61, 70, 58, 30, -10, -4, -3, -3, 16, -17, -1, -10, -14, -12, 2, 15, -19, -15, -18, 18, 7, 8, -9, 27, 2, -8, -4, 31, 10, 8, -15, -13, 5, -27, -18, 12, 20, -7, -4, 15, -11, -9, -10, 5, -13, 2, -4, 3, 14, 2, 9, 47, 5, -28, -20, -9, 25, 37, 1, -9, -40, -31, -6, -29, -21, -12, -10, 2, -16, 0, 10, 0, -19, -18, -7, 9, -2, -35, -8, -48, -33, -64, -63, -26, -15, 17, -11, -3, -21, -12, -31, -22, -15, 16, 0, 9, -20, -9, 7, 2, -2, 7, 14, -13, -3, 9, -21, -41, -41, -35, -34, -1, 6, 2, -17, -8, -16, 11, -33, 2, 6, 39, 16, -1, -13, 1, 11, 1, 5, -12, 4, -5, 23, 19, -23, -18, -3, -21, -24, 13, 29, 12, -7, 10, -4, -23, -3, -20, 15, 24, 28, -7, -14, 10, 16, -2, 12, -14, 19, 12, 35, 0, 14, -4, -49, -21, 30, 17, 5, 30, 25, 23, -1, -21, -20, -25, -6, -5, 12, 14, -4, 11, -1, -17, 1, -6, -8, 36, 59, 1, 11, -56, -58, -31, 28, 30, 42, 45, 20, 24, 31, -2, 15, 31, 5, 16, 32, 6, 8, -13, -6, -5, 15, 0, -1, 77, 51, 9, -15, -34, -55, -61, 11, 8, 27, 23, 29, -23, -10, -4, -4, 46, 25, 26, -17, 36, 37, -6, 8, 19, 19, -6, -11, 74, 26, -24, -18, -28, -28, -66, 23, 27, 48, 31, 37, 3, -4, 14, 15, 29, 4, 38, 34, 53, 44, -16, -1, -12, 13, -18, 23, 65, 39, 0, 9, 16, -30, -48, 48, 64, 20, 22, 16, 6, -14, 10, -15, -44, -42, -3, 28, 19, 48, -18, 8, 2, 6, -29, 39, 68, 27, 4, 20, 22, -10, -36, 57, 46, 23, 11, -4, 9, -49, -27, -39, -79, -46, -22, 0, 24, 33, -20, -3, 15, -14, -35, 21, 3, 41, 39, 25, 18, -1, -52, 31, 50, 20, 43, 27, -9, -32, -58, -75, -59, -40, -69, 9, 8, 30, 3, -14, 0, -6, -12, -7, -2, 4, 1, -22, 4, -32, -26, 34, 31, 28, 48, 19, -22, -69, -51, -29, -59, -41, -25, -3, 7, 14, -3, -3, -17, 6, 9, 38, 9, 13, -14, 5, -28, -26, -14, 6, 30, 41, 17, -2, -18, -56, -56, -45, -98, -65, -29, -9, 13, 14, -20, -1, 16, 5, 31, -25, -21, 8, -28, -19, -34, -31, -8, 38, 20, 17, 35, 38, -13, -49, -71, -98, -90, -52, -18, 4, 7, 17, -14, -18, 7, -12, 43, -41, -46, -57, -59, -31, -46, -36, 4, 16, 37, 2, 47, 44, -7, -64, -72, -64, -62, -57, -16, -9, -2, 1, 10, -17, 13, 6, 61, 11, -22, -72, -52, -43, -49, -36, -14, 43, 32, 6, 18, 44, -4, -28, -22, -17, -45, -68, -46, -27, -15, 18, -12, 1, -2, 14, 42, 34, 1, -29, -35, -22, -42, -39, -27, 8, 10, 35, 19, 20, -17, -70, -84, -60, -101, -99, -41, -51, 3, -15, 17, 15, 11, -13, 57, 55, -6, -43, -36, -30, -37, -38, -31, 10, 9, 18, 22, 29, 18, -42, -70, -83, -55, -35, -55, -7, -36, -22, 13, -13, 2, 5, 73, 27, -64, -37, -28, -49, -38, -54, -35, -29, 19, 19, -1, 10, 25, -57, -45, -43, -67, -43, -47, -44, -12, 3, 10, 1, -17, -19, 43, -9, -37, -67, -63, -39, -23, -5, -20, -15, 2, -5, 10, 12, 4, -35, -40, -27, -50, -31, -23, -8, -32, -12, -7, 11, -3, 3, 13, 26, -32, -18, -39, -39, -42, 9, -22, -35, 63, 1, -4, 5, -7, -50, -27, -39, -36, -41, -13, -14, 3, -5, 14, -20, 19, -10, 1, 5, -26, -15, -31, -32, -38, -4, 0, 26, 22, 7, -21, 11, -37, -42, -31, 22, -45, -3, -8, 8, 7, 26, 9, -14, 3, 9, 34, 13, -6, 1, -13, -21, -33, -53, -10, 12, 50, -42, -7, -3, -39, -10, -26, 5, -28, -30, -4, 10, -8, 5, -6, 13, 9, 9, -12, 11, -1, -23, -7, -25, -3, -25, 8, 2, 19, 5, 1, -18, -29, -26, -12, 22, -29, -26, -11, 5, 9, -5, 16, -11, -17, 7, 9, -12, 0, -11, -38, -21, -25, -6, -3, 43, 2, 21, 10, 9, -14, -18, -10, 14, -1, -17, 2, -9, 8, 15),
  115 => (1, -15, 10, 4, -7, -3, 9, 14, 4, 1, 15, -4, -10, 2, 9, 22, -34, 9, -26, -15, 2, -2, 20, 12, 8, -3, 10, -10, 1, -3, 5, -14, -7, -15, 10, -2, 12, -10, -4, -13, 30, 48, -17, -42, -18, -27, -29, 16, 79, 12, 10, 9, 8, -13, 17, -2, 10, 0, -2, -17, -3, 10, -10, 5, -7, -13, 34, 9, 12, -29, -57, -81, -37, 4, 25, 91, 116, 48, 33, -4, -11, -15, -6, 16, 12, 15, -10, -19, 3, 10, 5, 3, 7, 54, 36, 34, 9, -2, -17, -29, 0, 18, 19, 32, 18, 20, 21, 19, 9, -18, -10, 20, -7, 16, -11, 7, -17, 8, -5, 17, 54, 71, 50, 9, 12, -11, -27, -13, 10, 31, 46, 37, -12, 16, -3, -6, -24, 3, 3, -4, -19, 11, 20, -8, -13, 13, -2, 46, -5, -38, -40, -28, -18, -23, 14, 39, 36, 10, 21, 25, 6, -10, -28, -10, -4, -18, 4, -13, 8, 12, -8, 12, -4, 7, -6, 14, -69, -46, -4, -14, -25, -4, 43, 50, 38, -1, 21, 17, -24, -37, 7, -25, 6, -10, -1, -13, -6, -11, 7, -1, 0, -10, -4, -22, -37, -3, 7, -28, -15, -10, 33, 20, -6, -13, 46, -3, -31, -49, -47, -13, -21, -32, 5, -21, 17, -19, -17, -20, -2, 2, -20, -31, -23, 40, 17, -27, -44, 10, 23, 12, 22, -6, -1, -20, -34, -56, -71, -22, -29, 0, -21, 1, -14, 8, -15, -1, 3, -10, -68, -32, 3, 31, -14, -61, -14, 12, 9, 34, -8, 10, -21, -32, -19, -37, -58, -41, -39, -21, -3, -3, 14, 8, -2, -4, -5, -37, -36, -22, -22, -1, -21, -69, 0, 23, 45, 32, 30, 3, -11, -24, -31, -37, -63, -47, -44, -4, -23, 6, 15, -18, 3, 8, 6, -19, -31, -24, -5, -27, -73, -28, 4, 36, 17, 14, 34, 1, -48, -22, -26, -57, -66, -43, -65, -37, 12, -19, -10, 7, -1, 7, 6, -12, -22, 3, -58, -11, -46, -23, 0, 30, 45, 22, 16, -7, -55, -61, -1, -6, -53, -58, -24, -49, -2, -24, -19, 18, -2, 19, -7, -58, -12, -15, -49, -33, -27, 4, 35, 52, 14, 47, 13, -44, -40, -66, -7, 4, -13, -49, -26, -3, 4, 11, -4, 12, -1, 11, -12, -30, 11, -72, -71, -55, -52, 6, 13, 13, 36, 24, 8, -57, -29, -42, -46, -11, -17, -1, -9, -19, 1, -3, 15, 15, 7, 20, -10, -31, -11, -53, -93, -67, -56, 31, 34, 24, 28, 39, -13, -51, -4, -14, -13, -3, -5, 19, 17, -41, -8, 7, -3, -9, -3, -3, -32, -28, -41, -75, -71, -87, -27, 43, 4, 23, 29, 4, -17, -27, 3, 1, -31, -14, -20, 3, 10, -21, -9, -1, 11, 13, 2, 0, -3, -48, -81, -89, -86, -61, -28, 54, 27, 26, 6, 4, -16, -3, 8, -11, -2, 19, 10, 2, -17, -18, -2, -25, -18, 13, -10, -5, 14, -47, -54, -66, -62, -49, -4, 55, 18, 28, 19, 2, -17, 12, 10, -16, 7, -16, -33, -33, -26, -1, 5, 3, 2, -10, 2, 6, 23, -26, -37, -36, -69, -44, 40, 56, 46, 26, 60, -2, -39, -24, -8, -29, -14, -33, -50, -52, -24, 0, 9, 13, 15, 3, -1, 8, -15, -22, -5, 8, -26, -26, 31, 48, 29, 63, 70, 16, -30, -55, -32, -31, -16, -28, -22, -32, -19, -35, 18, -17, 10, 3, 18, -2, -66, -48, 11, -26, -41, -32, 25, 45, 23, 12, 2, -25, 5, -33, -25, -57, 13, 3, -13, -25, -17, -1, -10, 5, -16, -14, -18, 14, -30, -61, -2, -37, -32, -12, 29, 7, -2, 6, 19, 3, -18, -39, -12, -38, 3, 5, -42, -65, -21, -16, -27, -12, 3, 3, 14, -11, -12, -59, -42, -21, -24, -20, 42, 20, 10, 21, 31, 35, -25, -35, -34, -8, -6, -7, -23, -13, 1, 37, 21, -8, -15, 7, 0, 20, -11, 6, -38, -31, -30, -11, 31, 18, 27, 32, -16, -12, -22, -41, -47, -37, -4, 42, -38, -12, -13, 26, 12, 5, 5, 13, -19, 7, -11, 2, -2, -12, -34, -2, 11, 12, 11, -6, -25, -49, -20, -37, -35, 7, 16, -20, 11, 21, -2, -23, -13, -7, 7, 14, 6, -5, 5, -18, -25, 8, -23, -2, 24, 32, 31, 0, -21, -35, -34, -56, -26, -31, -27, -17, -22, 41, 9, -18, 14, -24, -18, 9, -9, 8, -17, 11, -11, -10, -7, 29, 6, 16, 19, 33, -22, -40, -46, -81, -52, -28, -19, 25, -20, -14, 9, 4, -3, 20),
  116 => (12, -15, -9, 10, -6, -19, -17, -1, 4, 9, 2, 15, -7, -15, 17, -27, -16, -26, -2, -11, -3, 15, 3, -14, -6, 4, 4, -7, 21, -18, 7, 13, -1, 12, -7, -17, -11, -1, 1, 17, 28, -2, -4, -19, -30, -21, 2, -2, 12, 17, -8, 9, -8, 7, -19, -7, -9, -12, -15, -16, -16, -4, 14, 14, 20, 14, -7, -31, -32, -8, -22, -32, -49, -1, -9, -15, -2, 9, -12, 4, -7, -16, -17, -2, 2, -2, -11, -6, -18, -2, -8, -12, 22, -40, -42, 8, 21, 21, -18, -22, -29, -29, -31, -2, -3, -8, 1, 16, -16, -12, -14, 6, -12, 12, -5, 9, -3, 8, -15, -19, -43, -14, 12, 20, 33, 7, -10, -8, -16, -28, -37, -36, -41, 9, -14, 4, -21, 7, 5, 12, -18, 18, -2, -16, -12, -18, -11, -45, 4, 1, 21, -8, -5, 5, 2, 10, 8, -15, -35, -63, 0, 9, 7, -14, -1, 2, -3, 12, 20, -19, 17, -5, -18, -17, -18, 4, 12, 9, -5, -28, 39, 34, 23, 6, 9, -8, -10, -31, -44, -45, 13, -14, 19, -20, -13, -15, -8, -9, 7, -18, 12, 3, 14, 22, 17, -30, -20, -31, 7, 19, -16, -8, -8, -21, -32, -43, -5, -41, -12, 26, -14, 11, -16, -5, 0, -3, -19, -10, 17, -13, 5, -3, 27, 22, -16, -61, -21, -32, 5, -3, -18, -6, -5, -31, 1, -19, 2, 11, -13, 13, 3, -2, 15, 13, 18, -10, 18, -5, 22, 43, 52, 24, -19, -1, -49, -49, -18, -33, -41, -29, -52, -19, -25, -12, -33, -6, 27, -3, -15, 15, -2, 3, 18, -2, -11, -9, -23, 2, 2, 19, -1, -16, -54, -52, -37, -39, -46, -30, -42, -6, -23, 18, -2, -43, 2, -20, -2, 13, 0, 20, 2, -13, -11, -17, -27, -3, 12, 11, -22, -3, -35, -68, -84, -90, -87, -59, -31, -28, -22, -13, -14, -63, -26, -7, -16, -8, 14, -15, -9, -7, 25, -8, -5, -14, 16, -3, 4, 36, 47, -11, -21, -71, -90, -77, -73, -82, -27, -65, -28, -83, -54, -13, 12, -20, -14, -16, -4, -6, -31, 24, 0, 14, -6, 6, 7, 32, 10, 41, 24, -4, -27, -40, -94, -55, -64, -44, -47, -57, -84, -12, -5, 11, -8, 12, 1, -2, -20, 43, 47, -3, -29, -36, 11, -16, -21, -6, 13, -2, -5, 11, -17, -61, -40, -53, -39, -86, -60, -56, 21, 2, -1, -18, 11, 2, -12, 37, 60, 17, -22, 3, -10, -21, 6, 1, 12, -14, -2, 8, -15, -27, -26, -37, -56, -78, -49, -42, -17, 2, 15, 7, -18, 2, 8, 10, 10, 10, -1, -8, 11, -4, 22, 10, 39, 23, 15, 6, 13, 14, -14, 11, 13, -28, -67, -54, -24, 0, -10, -16, -16, 11, 16, -19, 1, -7, -18, -17, -12, 27, 28, 9, 25, 29, 31, 11, 18, 59, -15, 20, 18, -19, -33, -14, -20, 23, 3, -13, 0, 11, 32, 34, 20, -6, -7, 10, 22, 37, 9, 12, 21, 33, 13, 52, 39, 33, 9, 14, 14, -9, -13, 9, 4, 10, -3, 8, 5, 5, 45, 20, -10, 14, 30, 9, 17, 41, 49, 52, 63, 40, 33, 56, 39, 30, 13, 14, 22, 19, 4, -8, 62, 21, 0, -6, -20, -14, 8, -51, -22, -6, 20, 23, 10, 19, 46, 29, 64, 57, 56, 30, 70, 40, 23, 49, 31, 7, 28, 5, 21, 28, -19, -16, -19, -3, -6, -45, -48, 4, 1, 20, 3, 10, 23, 26, 34, 57, 66, 88, 45, 50, 70, 54, 67, 65, 45, 4, 22, 7, 4, 14, -4, 6, -40, -77, -64, -10, 43, 2, 4, 10, 24, 1, 35, 43, 62, 69, 75, 59, 35, 47, 50, 58, 77, -1, -9, -20, 7, 15, -18, 11, -37, -35, -65, -18, 12, 4, -11, 17, -22, 2, 15, 37, 11, 16, 42, 41, 21, 52, 68, 59, 63, 54, 7, -27, 20, 10, 17, 20, 47, -24, -27, 0, -2, 13, 14, 17, -6, -3, -16, 25, 16, 17, 33, 25, 36, 68, 62, 58, 70, 33, 30, 21, -15, -19, 7, -15, 20, -9, -18, -3, 51, 2, 3, -12, 3, 4, 21, 10, 24, 15, -3, -16, 16, 46, 53, 39, 58, 66, 41, 55, -3, 0, 15, 10, -9, 7, -26, 10, 1, 3, 21, -8, -8, -41, 10, -23, 7, 22, 3, -2, 3, 36, 38, -12, 20, 72, 47, 57, -18, 10, 7, 12, -1, 0, 34, 43, 19, -1, -24, -12, -18, 0, -31, -48, -22, 4, 46, 24, 43, 8, -4, 13, 9, 23, 10, 38),
  117 => (14, -1, 17, -11, -2, 7, 19, -18, 8, 4, -4, -20, -1, -17, 7, -4, -52, -17, -29, -48, -16, -3, 6, -6, -1, -3, -13, -1, 8, 1, -8, 15, 4, -3, 6, 10, -1, -9, -14, -11, -47, -44, 0, -12, -10, -14, -20, -13, -41, -4, -12, 17, 13, -8, -2, 1, -13, 5, -21, -9, 16, -3, -15, 15, 20, -17, -39, -22, 2, -5, 7, 12, 31, 40, 3, 23, 3, -4, -5, 28, -13, 22, -15, 3, 18, 0, -1, -5, 8, -4, 12, 2, -2, -16, -13, -23, 20, 43, 25, -13, -30, -29, -5, -4, 2, 35, 27, 30, -1, 4, -10, 7, 15, 18, 8, -2, -1, 8, -2, -28, -6, -18, -28, 41, 59, 14, -11, -18, 14, -17, 30, 22, -1, 22, 7, 24, -4, -11, -4, -6, -13, -5, -17, 18, 9, 17, -18, 1, -29, -53, -3, 63, 57, 15, -23, -11, 16, 24, 20, 9, -8, 9, 8, 33, -1, 29, 8, -10, -19, 12, 1, 18, -17, -3, 0, 10, -34, -12, 39, 49, 57, 1, 6, -57, -28, -3, 1, 24, -4, -6, 29, 17, -31, 0, -6, -4, -10, -14, 16, -3, 3, -7, -11, -22, 35, -2, 40, 31, -12, 17, -21, -34, -14, -14, -24, -29, 2, -2, -31, -5, -24, 27, -17, -1, -11, -3, 15, 2, -6, 4, 15, 31, 6, 23, 27, 28, 12, -4, -35, -18, -40, -13, -37, -67, -27, -63, -32, -36, 21, -10, -6, -5, -5, -13, 1, 1, -7, -17, -17, 4, -2, -16, 26, 19, -4, 0, -22, -48, -58, -23, -10, -70, -61, -43, -57, -40, 9, 11, -15, -18, -13, -10, 13, 16, -20, -19, -47, -8, -38, -10, 24, -6, -6, -29, -35, -80, -53, -63, -88, -86, -75, -86, -53, -42, -29, -7, -45, 13, 19, 17, -21, 8, 8, -39, -68, -47, -9, 13, -3, -5, -11, -8, -49, -33, -79, -59, -51, -55, -54, -22, -33, -44, -32, -18, -26, 17, -2, 15, -7, -15, -20, -24, -99, -54, -36, 7, -17, -30, -42, -22, -7, -8, -12, -13, -31, -17, -31, -25, -26, -51, -52, -62, -36, -2, -12, 18, -9, -5, 27, -21, -68, -42, -67, -24, -42, -45, -8, -32, -39, -9, 28, 12, 1, 34, 2, 2, -8, 6, 15, -45, -18, -47, 12, 10, 13, 2, 0, 32, -19, 10, -18, -25, -16, -10, 23, 13, 4, 18, 1, 38, 34, 36, 66, 65, 41, 24, -2, 13, 14, 23, -9, 11, 5, 11, -10, 53, 7, 34, -11, 16, 37, 48, 23, 26, 34, 16, 61, 51, 24, 43, 72, 80, 52, 8, 30, 3, 3, 9, 0, -7, -18, 16, 32, 51, 28, 19, 34, 55, 45, 44, 27, 3, 23, 47, 71, 25, 41, 29, 52, 70, 42, 20, 26, 23, 20, 14, 15, -12, 20, 6, 3, 49, 7, 29, 6, 25, 47, 47, 20, 7, 22, 39, 67, 47, 47, 41, 13, 11, 12, 20, 14, 28, 10, 29, -4, -20, -3, -11, 52, 43, 35, 3, 35, -2, 55, 39, 45, 23, 39, 41, 17, 33, 59, 23, 38, 14, 29, 1, 9, 24, 21, -1, -11, -20, 11, 6, 84, 36, -26, 9, 23, 24, 31, 44, 49, 28, 64, 17, 30, 57, 26, 12, 19, 11, 29, 21, -13, 45, 42, 13, -14, -5, -9, -15, 34, 46, 23, -7, 34, 18, 30, -3, 16, 21, 47, 73, 42, -15, 6, 7, 12, 20, 19, 39, 16, 5, 42, 52, 0, -16, 18, -18, 36, 31, -7, 25, -5, 8, -28, -2, 4, 23, 14, 14, 19, -6, 18, 2, 3, 29, 30, 14, -30, -17, -43, 14, 0, -9, 19, 6, 44, 25, -26, 20, 36, -29, -36, -34, -17, -41, -12, -39, -29, -30, 18, -17, -32, -41, -29, -5, -15, -14, -32, -6, -5, -12, 19, 20, 60, -23, -36, 7, 39, 17, -23, -20, -55, 10, -24, -40, -36, -45, -34, -61, -38, -41, -42, -57, -64, -18, -39, 12, -2, 13, 20, 20, 14, -9, -13, -1, -10, -46, -21, -6, -25, -1, -51, -28, -32, -82, -24, -60, -41, -67, -26, -53, -61, -57, -17, 14, -12, -4, 19, -17, 1, -24, 3, 16, 4, -18, -24, -47, -18, -13, -34, -12, -50, -66, -25, -35, -31, -32, -35, -45, -52, -57, -54, 15, -18, 15, 4, -7, 11, 62, -15, 15, -1, -22, -4, 0, -18, -25, -16, -31, 11, -32, -47, -27, -16, -30, -47, -17, -30, -13, -37, -41, -5, 14, 6, -20, 17, 23, 45, 73, 49, 46, 0, 5, 7, -8, -31, -12, 6, 14, -15, -39, -26, -23, 0, -12, 15, 21, -18, -19),
  118 => (18, 1, -3, -10, -8, -2, -11, 3, -5, 3, -7, -13, -7, 3, 13, 9, 3, -20, -35, 8, 17, 39, 16, 6, -9, 8, 2, -13, 17, -8, 18, -2, -7, -9, 14, -3, -15, 7, 15, 20, 12, 39, 21, -9, -36, -33, -15, -16, 9, 7, -10, -15, -16, 5, -2, 4, 19, -11, -18, -15, 16, 4, -3, 2, -9, 25, 29, 31, 15, 18, -33, -33, -51, -43, -15, -11, 24, 10, 14, -25, 10, -13, -6, -7, 6, 15, 5, -14, -4, -15, -14, 1, 10, 15, 16, -27, -39, -42, -57, -41, -44, -38, -67, -61, 17, 53, 12, 27, 31, 18, -12, -18, 2, 12, 12, 10, 2, -6, 7, 40, 16, -1, -42, -62, -72, -100, -65, -44, -55, -24, -20, 4, 52, 7, 17, 21, 28, -45, 19, 14, -4, -9, 6, -8, 19, 3, 0, -26, 8, 7, -28, -71, -59, -77, -49, -39, -47, -9, -5, 10, 23, 39, 67, 30, 0, 26, 14, -7, -18, 15, 6, 13, -4, 18, -34, -5, -13, 2, -30, -54, -31, -50, -62, -18, -42, 0, 14, 20, 44, 8, 72, 32, -15, -21, -28, -4, 17, -10, -13, -7, 3, 5, -3, -16, 7, -35, -67, -64, -40, -64, -43, -54, -6, -7, -13, 0, 38, 13, 29, 21, -34, -20, 2, 33, -15, -8, -7, 4, 3, -6, -4, -21, -57, -21, -55, -12, 21, -14, -4, -2, 29, 53, 65, 68, 80, 89, 45, 77, 46, 31, 58, 24, -8, 20, 7, 19, -10, -19, -15, -38, -25, -12, -14, 48, 24, 41, 11, 30, 29, 20, 39, 45, 54, 67, 28, 65, 65, 18, 38, 38, -3, 1, -20, -7, 6, 1, 63, -20, 1, 18, 12, 13, 18, 48, 28, 42, 20, 1, 41, 24, -16, 24, 10, 7, 18, 2, 33, 36, -14, -18, -6, -10, -13, 68, 65, 38, 81, 39, 31, 35, 26, 26, 6, 0, 46, 1, 36, 49, -6, 8, 8, 19, 33, -6, 7, 9, -9, 3, -17, 14, -38, 40, 47, 16, 61, 5, 1, 17, 15, 46, 35, 12, 24, -5, 21, 8, -56, -5, -5, -34, -19, -32, 13, 36, 17, 6, 16, -7, -28, 24, -24, 35, 34, 52, 40, 50, 32, 22, 51, 45, 17, 7, -23, 2, -35, 2, 4, -33, -17, 3, -36, 20, -11, 20, 4, -7, -20, 29, 46, 11, 29, 33, 2, 34, -24, 10, 24, 1, 7, -13, -33, 7, -8, -16, 10, -48, 8, 23, -20, 52, -6, -17, -1, -15, 3, 33, 34, -5, 2, 38, -8, -55, -11, -33, -17, -18, -8, -17, -17, -3, 21, -14, -15, -24, 5, 4, -28, 42, 6, 17, -11, 13, -1, 18, 52, 24, 27, 15, -40, -44, -25, -20, -2, -7, -11, -30, -26, -26, 2, -33, -53, -24, -32, 3, -20, 36, 18, -16, 16, -3, -7, 1, -4, -21, 19, -28, -31, -35, -22, 0, 2, 2, 23, -9, -73, -41, -28, -22, -14, -38, -36, 2, 34, -18, 18, 9, 5, -7, 19, -15, -4, -41, -35, -55, -60, -37, -17, -7, -15, -12, -9, -18, -56, -58, -25, -32, -25, -17, -8, 16, 43, 31, 9, -4, -19, 1, 2, 10, -16, -3, -31, -66, -17, 2, -7, 18, 18, 11, 24, -12, -63, -55, -46, -59, -3, 17, -38, 55, 82, 68, -5, 2, -6, -19, -2, 11, 8, 11, -19, -6, 4, -26, -2, 74, 9, 75, 26, -6, -39, -25, -37, -41, -17, -3, -16, 14, 75, 86, -2, -7, -1, 7, 49, 13, -19, -18, -11, -15, 30, 3, -6, 43, 23, 66, 8, -29, -23, 1, -25, -8, -8, 24, 7, 14, 29, 31, -12, -17, 3, -15, 6, -14, -23, -3, 14, -40, 6, 33, 33, 21, 30, 13, -12, -64, -73, -60, -1, 1, 27, 43, 58, 41, -5, 25, -9, -2, 8, -14, -9, -21, 5, 7, 2, -20, 24, 31, 47, 38, 38, 15, -17, -65, -48, -61, -63, -52, 10, 45, 60, 14, -21, 16, -14, 7, -12, -13, -20, -50, -19, -32, -27, 4, 31, 19, -6, 37, 34, 1, -29, -75, -87, -90, -38, -26, -21, 25, 26, 1, -17, 46, 13, 6, 11, 14, 27, 5, -10, 0, -8, -27, 1, 21, 42, 63, 7, -36, -37, -42, -90, -36, -4, -11, -21, 25, 52, 4, 2, 20, -17, -11, 3, 17, 5, 20, -27, -22, -21, 30, 17, -13, 20, 64, 36, -10, -39, -82, -85, -24, -9, 27, -16, -3, 0, -3, 8, 31, 13, -8, 7, 7, -19, -8, 20, 15, 17, 18, 38, 11, 8, -11, -31, -5, -19, -44, -44, -61, -37, -3, 28, -7, 23, 19, 24, 7),
  119 => (-10, 16, -11, 5, -17, 3, -1, 0, 2, 17, 2, -8, -5, -16, -5, -37, -14, -46, -11, -7, 15, -13, -19, -2, -14, 4, -19, 6, 8, 18, -3, 8, -16, 11, -3, 17, -10, -5, 12, 3, 7, -20, -35, -26, -12, -41, 0, -27, -2, -7, -20, -2, 3, 11, -17, 7, -3, 19, 7, 8, -21, -7, -2, 0, -12, 11, 27, 36, 9, -7, -32, -13, -27, -43, -60, -20, -2, 13, 23, 13, -11, -20, -2, 19, 11, -18, -17, 2, 16, 17, 12, 12, 13, 3, -24, -27, -50, -52, -45, -24, -22, -3, -4, 6, -9, -7, -6, 10, 0, 1, 3, 12, 15, 11, -7, -12, -13, -18, 5, 11, 32, -5, -62, -37, -52, -26, -49, 5, 12, 30, 13, -15, -83, -65, -21, -9, 17, -6, 8, -4, 19, 0, 11, -3, 9, 19, -15, -18, -10, -49, -30, -56, -54, -19, -11, 24, 29, 18, -7, -26, 5, -26, -20, -31, -12, 12, 19, 1, -8, -8, 18, -5, 9, 20, -4, -11, 9, 5, -21, -32, -70, -49, -32, 1, 21, 19, 25, -19, -17, -36, -51, -41, -19, 4, -8, -3, 6, -4, -20, -20, -5, -17, -1, 16, 26, 17, 4, -36, -24, -6, -21, -5, 6, 2, 10, 18, 27, 7, 13, -45, -17, 12, 28, 20, -1, 4, 10, -12, -11, -15, 18, 26, 27, 24, 31, -20, -31, -14, -20, -10, -25, -42, -32, -18, 11, 12, 42, -23, -49, 12, 26, -4, 0, -16, -3, 6, -9, -1, 21, 22, 22, 24, -6, -11, 31, 32, 48, 9, 2, -16, -10, -19, -34, -1, -1, 14, -2, -25, -16, 24, -17, 11, -17, -13, 13, -48, 7, 33, -15, -25, 0, -12, -1, 47, 38, -4, -19, -10, -6, -20, -5, -22, -29, -9, -15, -43, 9, 30, 12, 16, -7, 13, -20, -12, -4, 7, -6, 5, 1, -4, -10, -39, 0, -15, -40, -78, -31, -70, -78, -50, -60, -64, -52, -35, 13, 26, -15, -1, -9, -17, -6, -19, 16, -17, 8, 34, 37, 33, 27, 18, 54, 30, -17, -11, -39, -86, -56, -53, -108, -77, -39, -60, 3, 6, -8, -18, 8, -6, -15, 0, 17, -24, -14, -22, 36, -3, 24, 30, 32, 44, 31, 12, 9, -4, -4, -25, -93, -94, -42, -40, 7, 7, -8, -14, 14, 16, 12, 3, -20, -33, -86, -49, -24, -9, -11, 10, 50, 62, 13, 36, 19, 24, 6, -15, -20, -54, -42, -60, -16, 10, -10, 7, 5, 0, -10, -9, -9, -66, -70, -75, -63, -71, -69, -62, 1, 2, 7, 9, 26, 30, 14, -4, -4, -14, -17, -14, 4, 17, -9, 2, -4, 17, -23, -12, -22, -29, -30, -37, -37, -59, -52, -61, -33, -25, -34, -22, -35, 32, 43, 21, -7, -19, 32, -17, -6, -15, 15, -5, 3, 20, -22, 2, 2, -27, -19, -13, -9, -26, 8, -4, -8, -9, -15, -37, -44, -20, 33, 44, 26, -1, 30, 53, 0, -5, 4, 11, -3, -8, 23, 38, -7, 32, 29, 57, 25, 16, 13, 42, 32, 48, 16, 40, 0, -58, -48, 2, 28, 25, 52, 31, 55, 2, -5, -14, -15, -3, 50, 37, 43, 52, 39, 39, 19, -5, 16, 8, 51, 16, 23, 12, 0, -38, -27, -5, 4, 19, 51, 58, 65, -21, 0, -10, 4, 3, 60, 27, 65, 13, 27, 4, 6, -8, -10, 7, 10, 16, -4, 5, -2, 4, 16, 6, 5, 2, 14, 32, 41, -37, -3, -3, -15, -9, 32, 23, -10, -36, -67, -54, -65, -73, 4, -20, -7, -7, -6, -13, -21, -5, -25, -21, -5, -31, -41, -7, 34, -57, 13, 7, 1, 2, 21, 14, -30, -42, -45, -59, -43, -73, -26, -3, -30, -20, -19, -27, -9, -16, -5, -16, -4, -13, 8, 15, 39, -23, -16, -10, -10, -12, 8, 10, -22, -29, -13, -39, -68, -76, -76, -65, -62, -38, -41, -12, 19, -5, -4, -18, -8, -9, 4, 35, 30, -28, 1, -20, 8, 19, -16, 16, 7, -27, -12, -32, -67, -67, -57, -112, -70, -55, -34, -3, 10, 5, -7, 26, -28, 32, 21, -10, 6, -40, 8, -5, 3, -17, -17, 14, 5, 18, 36, 59, -11, -17, -29, 9, -7, 8, 14, 40, -11, -26, -19, -6, -32, 15, -27, -35, -52, -9, 14, -20, -18, -16, 2, -26, 7, 0, 34, 33, 26, 24, 31, 32, 54, 27, 19, 14, 43, 27, -2, -2, 7, 4, -31, -14, -12, 6, 11, 16, 17, -2, -2, 11, -10, 7, -24, 7, 21, -1, 25, 25, 18, 9, 23, 13, 12, 26, 42, 5, 12, -9, 8, -38, -6, -23),
  120 => (-13, -9, 16, 4, 18, -7, 12, -3, -6, -17, 16, 17, -1, 16, -16, -13, -38, -25, -23, -16, 5, -9, 28, 20, -14, 19, -4, 20, 4, 10, 14, 16, -14, 2, -4, 4, -15, 16, -18, 37, 1, 18, -1, -18, -81, -36, -53, -41, 6, -28, 6, 6, 3, 17, 3, -17, 1, 20, -13, 15, -5, -13, 16, 18, 0, 7, -15, 20, 0, -30, -28, -8, 23, 1, 35, -19, -6, -4, 36, 36, 29, -5, 3, 10, 12, 11, -17, -12, 7, -9, 18, -9, -19, 2, 35, 42, 25, -2, -34, -8, -43, -10, 12, 6, -26, -24, 21, -16, 3, -17, -10, -4, 15, 0, -7, -11, 10, 17, 11, 7, -40, 22, 23, 28, 29, -6, -27, -28, 5, 4, -2, -3, -1, -3, 8, -4, -20, -13, 5, 1, 14, 9, 15, 0, -10, -7, 16, -44, 13, 64, 33, 45, -6, -16, -33, -9, 18, 20, 1, 0, 21, 11, -7, -17, -30, -28, -3, 4, -16, 19, -7, -20, 17, -8, -30, 8, 28, 36, 39, -12, -4, -29, -2, 8, 2, -16, 20, 7, 13, -21, -25, -29, -11, -13, -2, -4, -2, -18, 17, -19, 14, 1, 34, 30, 5, 2, 1, -21, 7, 8, 31, 14, -8, -21, 8, 14, 6, -25, -34, -76, -39, -27, -49, -4, 13, 12, 9, 19, 0, -18, -2, 10, -35, -28, -68, -66, -16, 19, -1, 14, -12, -8, 7, 11, -6, -55, -74, -44, -42, -33, -18, -23, 0, -10, -7, 18, 21, -18, 5, -43, -87, -86, -106, -61, -52, 24, 28, 23, -11, -4, 30, -8, -40, -21, -9, -20, -31, -32, 3, -2, -6, 13, -20, 15, 17, 25, -44, -93, -104, -116, -110, -31, -20, 18, 37, 43, 3, 24, 33, 6, 18, -8, 12, -22, -5, 16, 20, 39, -7, -14, 13, -8, 20, -27, -113, -147, -107, -81, -72, -20, 5, 62, 24, 26, -10, 20, 38, 44, -3, -15, -28, 0, 32, 38, 37, 37, -9, -6, 3, -2, 6, -10, -88, -84, -51, 10, 0, -21, 40, 33, 8, 17, 35, 14, 26, -12, -27, -31, -21, -7, 9, 5, 24, 34, -10, 7, -18, 0, 34, 50, -13, -8, 15, 62, 13, 36, 33, 66, 39, 43, 58, 23, 4, 1, -2, -37, -22, 4, 1, -1, 2, 31, 6, 6, 10, 5, 50, 66, -10, 9, 22, 10, -22, 29, 59, 62, 47, 30, 15, -5, -4, 0, -33, -10, -35, -15, 6, -37, -5, -29, 0, 14, 6, -18, 26, 45, -35, 19, -18, -71, -3, 24, -5, 36, 67, 9, 16, 7, 14, -20, -30, 12, -19, -17, -18, -18, -21, -5, -2, 17, -16, -9, 56, 26, -20, -20, 8, -23, 49, 29, 9, 6, 4, -8, -13, -14, -47, -49, -30, -4, -70, -59, -26, -24, -1, 8, -12, 16, 14, 21, 73, 57, 16, 28, 18, 20, 59, 18, 12, 52, -11, -15, -35, -20, -47, -66, -46, -44, -79, -51, -23, -8, -16, 19, -6, -8, -20, 3, 28, 66, 8, 22, 13, 17, 58, 6, 51, 21, 3, 5, -47, -38, -41, -79, -66, -66, -82, -34, -39, -31, 2, 6, 9, 3, -18, 20, -12, 25, 30, 33, -11, 14, 25, 4, 42, 33, -3, 5, -9, -13, -9, -52, -48, -47, -90, -51, -47, 9, -19, -5, 18, 5, 20, 17, -30, -36, 21, 29, 10, 10, 45, 41, 27, 5, -30, -33, -5, -31, -33, -34, -37, -12, -7, 4, -39, 6, 5, 5, 8, 4, -17, -19, -11, 6, -9, 10, 18, 20, 75, 42, -18, 3, -10, -4, -4, -25, -47, -56, -57, 5, 18, 1, 1, 6, -10, 14, -5, 11, 11, -9, -11, -7, -6, 10, -1, 26, 55, 47, 12, 3, -22, -10, -37, -33, -82, -79, -98, -52, -57, -24, 27, 3, -1, -3, 0, 7, -12, -1, 21, 23, -47, 25, 9, -8, 12, 1, 30, -9, -29, 11, -30, -41, -36, -93, -35, -23, -35, -54, -15, -9, 1, -15, -8, 7, -2, 7, 81, 95, -6, -13, -23, -10, -22, -4, -13, -9, -19, 3, -11, -41, -18, -20, -8, -29, -23, -29, -40, -24, -2, 21, -1, 14, 21, 5, 40, 38, 3, -12, -43, -43, -54, -79, -37, -49, -43, 8, -30, -41, -25, -48, -25, -11, -40, -18, -24, -13, 35, -11, -1, -11, 19, -13, 28, 24, -36, -24, -30, -74, -28, -43, -35, 1, -7, -29, -46, -8, -42, -13, -30, -26, 4, -1, 1, 4, 21, 10, 13, 5, 16, 8, 12, 2, -20, -15, 8, 14, -27, -38, -3, -15, 8, -4, -53, -26, -52, -49, -29, -17, -21, 3, -19, 2, -27, 13),
  121 => (-14, 6, -1, -7, 17, -20, -19, -20, -12, -20, 8, 18, -1, -14, -2, -1, -22, 14, -4, -7, -18, 0, -19, 15, 13, -6, -14, 1, 18, -11, -14, 6, 5, 8, 12, 19, -13, -15, -15, 3, 11, -19, 9, -40, -13, -12, -18, -8, 3, 6, -9, -14, -13, -4, -11, -1, 13, -19, 13, -6, -7, 5, -2, -7, 8, -8, 2, -1, 10, 8, -24, -25, -44, -21, -29, -16, -38, -6, 9, -18, -32, -5, 7, -19, -10, 1, 11, -8, -4, 3, -6, -14, 5, -18, -21, -5, 19, -37, -71, -111, -74, -70, -66, -60, -46, -40, -9, -19, -41, -39, 16, 7, -9, 8, 11, -15, 6, -5, -14, 13, -25, -21, 25, -21, -68, -83, -83, -129, -134, -111, -95, -62, -56, -53, -4, -4, 22, -21, 14, -18, -16, -19, 2, -19, 1, -6, -18, -22, -19, -51, -31, -75, -51, -1, -50, -114, -115, -107, -128, -122, -53, -57, -24, 13, -7, -8, 5, 18, 10, 12, -14, -12, 17, -1, -9, -29, -47, -24, -24, -54, -56, -65, -58, -34, -47, -35, -37, -5, -27, 6, 34, 58, -3, -6, -16, 6, -20, 6, -12, 19, -9, 7, -11, -72, -33, -37, 29, 36, 50, 30, 33, 7, 24, 25, 19, 24, 10, 20, 29, 49, 26, 3, -63, 1, -12, 2, 0, -12, 17, -4, -21, -24, -21, -4, 18, 19, 19, 28, 27, 4, 40, 15, 33, 38, -4, 27, 44, 52, 29, 36, -18, -17, 15, 10, 19, -15, 16, -7, -24, -11, -29, -42, -1, -3, -16, -14, 32, 14, 12, 23, 47, 64, 23, 24, 14, 8, -10, 44, -17, -20, -6, -18, -9, 14, -5, -8, -47, -10, -10, -46, -16, -40, -38, -29, -8, 12, -5, 25, 45, 80, 42, 16, 20, 1, 10, 23, 10, -26, 13, 14, -12, 14, 3, 7, -47, 12, -4, -24, -13, -22, -51, -63, -42, -21, -62, -44, 3, -13, -11, -31, -10, -60, -20, 5, 18, -17, -14, -19, 15, 10, 1, -4, 42, -1, 2, 23, 21, -15, 7, -15, -20, -41, -38, -45, -44, -52, -74, -47, -35, -61, -64, 28, 75, 44, -10, -4, 3, -5, -16, 82, 37, 57, 59, 63, 35, 65, 37, 15, -11, -3, -28, 4, -4, -22, -5, 2, -28, -31, -8, 22, 42, 30, -2, 10, 17, -12, 38, 83, 60, 48, 43, 34, 16, 22, 5, 37, -15, -6, 8, -15, 44, 7, -14, 2, -4, -23, 3, 1, 45, 25, -18, -19, -1, 2, 67, 59, 60, 18, 4, -13, 20, -28, -12, -1, 6, 10, 6, 26, 11, 9, -4, 9, -13, -3, -30, -34, 7, 53, 16, -9, 18, 9, 62, 58, 32, 7, -9, -16, 15, 12, 29, 40, 52, 26, 24, 37, 19, 46, 27, 7, 5, -4, -19, -12, 11, 81, -12, -13, -14, -11, 15, 53, -3, 22, -11, -30, -23, -15, -27, 0, 4, 2, -4, 15, 49, 13, 5, 12, -7, 19, 11, -15, -7, 64, 17, 9, 19, 0, -10, 16, -28, -62, -106, -73, -55, -38, -33, -60, -58, -36, -53, -39, 2, -21, -22, -18, -24, -7, -38, -70, -22, 42, 13, 7, -20, -1, -8, -19, -57, -72, -88, -112, -44, -1, -5, -30, -49, -25, -37, -47, -37, -12, -15, -9, -12, -28, -41, -47, -27, 32, -14, 9, 17, -3, -26, -54, -66, -59, -49, -62, -25, -9, 4, -17, -9, -37, -27, -43, -27, -44, -15, 20, -3, 32, 2, -14, -15, 39, 9, 16, 12, 10, -46, -42, -74, -55, -22, -33, -14, -3, 2, -23, -26, -3, -13, -6, -5, -38, -7, -11, -6, -24, 2, 11, 62, 49, 16, -12, 3, 1, 8, -8, -37, -42, -21, -43, -16, -9, 22, -29, 14, 10, 18, -40, -4, -21, 14, 29, 15, 23, 8, 37, 76, 14, 9, -18, 5, 18, 3, -23, -6, -35, -23, -3, 1, -5, 29, -18, 16, 13, -14, -33, -38, -2, -7, 2, 10, 7, 6, 24, 62, 42, 20, 13, 15, -9, 15, 5, -21, -5, -4, -38, -22, 5, -11, -20, 6, -20, -21, -11, -23, -31, -32, -8, 26, 15, 39, 57, 38, 29, -4, -6, 17, 15, 57, 40, 22, 40, 30, 1, 10, -9, -2, 20, -12, -7, -2, -30, -41, 2, -12, -4, -25, 5, 24, 57, 55, 26, 18, -2, -6, 13, 25, -4, 4, 32, 32, 20, -6, 13, 27, 24, 35, 54, 10, -42, -54, -34, -30, 13, 16, 22, 20, 31, 22, 8, -12, 3, -13, 0, -1, -10, 3, 35, 10, -4, 18, 49, 55, 48, 63, 37, 8, -8, -65, -46, -20, 16, 27, 30, 25, 25, 25, 11),
  122 => (-2, 15, 5, 16, 2, 13, 6, 9, -1, 5, -13, 1, -7, -11, 1, -48, -14, -26, -40, 1, 26, 62, 50, 12, -4, -15, 16, 11, -15, -7, 16, -15, 2, -13, 8, -16, 20, -17, -2, -11, 30, 28, 68, 67, 68, 66, 68, 54, 81, 27, 39, -20, -5, -19, -3, 10, 19, -12, -15, 10, 6, -19, -5, -6, 14, -11, 28, 51, 1, 50, 45, -3, 39, 28, -16, -2, 23, 60, 26, 12, 7, -17, -2, 17, -16, 8, -17, 14, -20, -19, 6, -2, 8, -34, -17, -31, 2, 18, 43, 27, 22, -28, -23, -19, -28, 14, 9, -20, -1, 12, -10, 16, 12, 2, -11, -1, 8, -12, 4, 2, -33, -24, -43, 24, 42, 49, 18, 9, -6, -9, 29, 16, 36, 14, -2, -23, -9, 30, -4, 20, -12, 11, -2, -12, 19, 0, -27, -45, -11, -28, -20, -4, -18, -21, 3, -3, -20, 7, -4, -4, 2, 3, -17, -36, -57, 5, -14, -6, 12, -12, 18, 12, 13, -15, -62, -11, 17, 12, -21, -21, -13, -7, -4, -12, -8, -27, -52, -12, -25, -43, -5, -53, -66, -8, -10, -5, -1, -3, 10, -18, 14, 19, -23, 9, 37, 39, 32, 12, 3, 1, -6, -23, -30, -19, -1, 0, -26, -30, -29, -33, -63, -48, 0, -12, -11, 10, -13, -16, 12, 12, -2, 37, 73, 87, 56, 64, -2, -21, -14, -24, -22, -37, -44, -9, -57, -55, -73, -73, -69, -35, 4, 23, 6, -17, 2, 11, 10, 16, 2, 63, 60, 45, 23, 22, 57, -10, -4, 1, -26, -25, -20, 3, 3, -31, -8, -46, -53, -16, 15, 36, 5, 5, -3, 2, -17, 13, 41, 85, 50, 54, -3, 9, 47, 30, 32, 4, -15, 4, -8, -4, 4, 24, 29, -24, -48, 12, 38, 59, -12, -15, 11, 14, 14, -6, 59, 58, 53, 37, 37, 14, 56, 47, 38, 30, 43, 12, 52, 13, 10, 8, -9, 1, 3, -11, 26, 45, -3, 13, -6, 19, 7, -22, 17, 40, 6, 3, -1, 13, 66, 19, 24, 72, 30, 29, 43, 28, 16, -5, 1, -17, 6, 10, 19, 15, -3, 2, -9, 5, -13, -35, -13, 27, -12, 3, 16, 17, 19, -2, 37, 55, 26, 18, 63, 29, 33, -3, 24, 23, 20, 9, 26, 22, 16, -13, 12, 13, -50, -10, 9, 21, 12, 0, 15, -17, -16, -9, 25, 26, 47, 24, 37, 34, 34, 26, 10, 31, 63, 7, 9, -11, -19, -7, -1, -7, 11, 4, -25, -7, -7, 16, 0, -15, -21, 5, 5, 9, 51, 12, 21, 18, 3, 32, 10, 4, 22, 65, 12, 11, -13, -19, 21, -16, 5, -36, -19, -16, -18, -22, -56, -52, -34, -44, -27, 19, 17, 22, 52, 13, 45, 35, 22, 37, 54, 56, 31, -13, 4, -17, -15, -7, -28, -25, -36, -41, -87, -48, -51, -24, -33, -20, -31, -23, -10, 9, 10, -2, 5, 11, 37, 61, 82, 56, 17, 30, 12, 14, 1, 5, -6, -21, -27, -55, -49, -63, -66, -58, -37, -33, -16, -21, -14, -7, -21, -31, -17, 7, 22, 48, 39, 32, 24, 17, 19, 3, -15, 2, 11, -34, -44, -42, -28, -27, -83, -38, -63, -31, -8, -42, -2, -4, 0, -34, -1, 23, -2, 8, 11, 18, 17, -19, -16, 9, 11, -17, -29, -56, -61, -20, -22, -17, -51, -69, -86, -60, 0, -44, -24, -21, -38, -38, -23, 9, 11, -19, 16, -6, -27, -2, 15, -15, -10, 8, -7, -36, -47, -35, -26, -47, -75, -59, -54, -68, -42, -37, -46, -61, -59, -38, -18, 8, -12, -23, -9, -9, -29, -32, 1, 2, -2, 7, -4, -10, -18, -40, -30, -55, -94, -89, -54, -39, -9, -28, -54, -91, -46, -37, -16, 35, -27, -38, -15, -16, -42, -57, 14, -9, 14, 19, 13, -22, -43, -38, 4, -39, -51, -35, -75, -25, -1, -46, -29, -87, -102, -58, -33, -19, -33, -37, -39, -36, -27, -16, 9, 14, 0, -10, -18, -46, -31, 14, -38, -44, -20, -24, -23, -35, -18, -33, -47, -68, -55, -61, -103, -73, -45, -13, 1, -42, -60, -40, -16, -3, 14, -17, 15, -5, 4, -53, -54, -51, -2, 10, -5, -13, -6, -17, -18, -20, -76, -61, -75, -62, -44, -13, 26, -29, -43, -11, 4, -18, 13, 14, 11, 7, -26, 9, -11, -10, 17, 19, -45, -17, -15, -24, 3, -21, -62, -56, -73, -77, -51, -31, 6, -25, -20, -3, 15, -1, -14, -3, 15, -7, 11, -5, -12, 5, -26, -13, -44, -59, -3, -49, 30, 3, 21, -9, -24, -30, -26, 5, 34, -1, 0, -6),
  123 => (-13, 19, 5, 12, -1, 16, 10, -17, -12, 14, 18, -20, 7, -13, -9, -10, 5, 9, -10, 15, 20, 17, 16, -12, 9, -6, 19, -12, 5, 12, 5, -1, -10, -6, 14, 19, -5, 7, -18, -19, -5, 6, -6, 3, -12, 0, 16, 7, -16, -6, 15, 20, 15, -13, -9, 12, -2, -17, -4, 5, 10, 7, 13, -12, -10, 13, 16, 10, -14, -16, -26, -36, -26, -22, -25, -23, -6, 10, 15, 26, 20, 2, -1, 15, 11, -10, -1, 17, -6, -3, 14, -1, 0, -2, 26, -8, -33, -49, -59, -25, -3, -5, -4, -19, -1, -19, 7, 1, 21, 8, 6, -2, 5, 9, -19, 11, -1, -5, 17, -8, 10, 9, 46, -37, -37, -14, -39, -31, -21, -21, -26, -18, -9, -11, 8, 12, -3, 18, 12, -18, 17, 10, 4, -16, -13, -15, -12, 12, 2, 39, 29, -8, -37, -2, -47, -6, -29, -49, -1, 4, 0, -22, 3, 57, 34, -2, -4, -1, -13, -9, -17, 10, -6, -9, 2, 19, 5, 43, -3, -8, -39, -83, -32, -35, -31, -34, 10, 14, -15, -9, 5, 16, 21, 21, -4, 6, 13, 11, -9, 15, -5, -17, -2, -3, 51, 40, 27, 16, -1, -24, -6, -10, 8, -7, 15, -24, -40, -17, -19, 12, 14, 38, -19, -12, 18, -10, -14, -4, -9, 12, -29, 22, 13, 38, 23, -27, 14, 12, -4, -25, -2, 5, 10, 0, -32, -14, -16, 6, 21, 27, -13, -2, -6, -14, 11, 2, 13, 15, -9, 21, -39, 1, -19, -57, -41, -53, -25, -45, -34, -23, -4, -15, -8, -7, -28, -9, -8, 23, -9, -7, -2, -2, 9, 17, -20, 19, -25, -9, -71, -86, -76, -75, -53, -46, -20, -50, -24, -37, -13, -50, -37, -25, -57, -6, -17, 15, 20, -23, 14, -11, 7, 7, -15, 18, -22, -33, -81, -63, -105, -103, -55, -52, -48, -25, -40, -22, -26, -25, -13, -33, -38, -20, -9, -26, -16, -3, -8, 10, 9, -16, -8, -24, -25, -53, -73, -65, -90, -81, -73, -64, -41, -45, -72, -40, -49, -49, -27, -34, -29, -24, -18, 0, 5, -24, -16, -15, -9, 15, -16, -1, -10, -35, -43, -37, -60, -45, -58, -42, -33, -31, -54, -41, -32, -35, 11, 0, -44, -28, 17, 12, 12, -2, -7, 18, 20, 11, -24, 22, 3, -16, -14, -19, -6, 8, -7, 18, 13, 5, 17, 38, 2, 35, 21, 9, 1, 16, 10, 29, 13, 71, 20, -5, -9, 3, 32, 55, 19, 31, 38, 10, 6, 33, 42, 15, 41, 53, 49, 29, 58, 53, 43, 40, 28, 3, 21, 29, 28, 62, 13, -3, 6, -16, 12, 52, 31, 50, 64, 57, 77, 84, 78, 82, 45, 35, 29, 59, 65, 38, 45, 37, 42, 48, 50, 23, 46, 38, 7, 8, -15, -13, 27, 40, 30, 54, 48, 38, 53, 55, 87, 51, 45, 27, 36, 3, 34, -2, 17, 41, 25, 10, 14, -2, 30, 54, -15, 20, -20, -18, 47, 53, 32, 33, 65, 7, 44, 57, 42, 69, 33, 27, 25, 5, -2, 13, -16, 10, 21, 2, 0, 10, -2, 41, 20, 14, -18, 9, 18, 42, 37, 4, -4, 2, 2, 23, 6, 34, 51, 32, 39, 0, -9, 19, -4, 5, -25, -10, -4, 24, -20, 17, -19, -10, 15, -16, 13, 29, 39, 7, -9, 11, 25, 29, 1, -5, 19, 25, 30, 0, -9, 15, -5, -10, 6, 4, -4, 3, -13, 15, 0, -13, 19, 20, -51, -47, -9, -8, -8, -16, 22, 57, -5, -1, 7, -11, 12, 1, -16, -13, -2, -18, -1, 2, 31, 26, -17, 11, 12, 7, 5, 5, -5, -50, -11, 14, 0, -2, 21, 39, 18, 30, -34, -7, -32, -18, -4, -35, -22, -22, -15, -13, -1, 21, -9, 23, 18, 5, 0, 2, -26, -29, 7, 9, -31, -5, 7, 36, 34, -1, -21, -8, 19, -13, -15, -24, -30, -28, -15, -32, -16, 3, -7, 1, -9, -5, 19, -18, -15, 15, 3, 44, 29, 33, 3, 18, 20, 21, 1, 28, 12, -15, -17, -3, -30, -20, 0, -28, -23, -11, 11, 26, -19, -11, 18, 7, -7, -25, 0, 13, 36, 50, 42, 25, 3, 11, 10, 25, 6, -11, -42, -23, 13, -3, -7, -33, -44, -10, 0, 9, 11, 0, -15, -16, -9, -12, -11, 22, 44, 0, -24, -13, 5, -29, -9, 23, -6, -51, -16, -4, -7, 2, -30, -46, -10, -17, -16, -5, 8, -15, 12, -15, -17, -12, 2, 11, 8, -1, -21, -39, -7, -6, -1, -32, 24, -8, -3, -8, -15, -32, -18, -5, -15, -17, -20, -25),
  124 => (11, -17, 15, 11, 0, -4, -20, -10, -14, -8, 8, 3, 7, -12, -9, -15, -10, -9, 13, 21, -11, -15, -9, -3, 13, 2, -13, 8, 4, 12, 20, 2, -21, 5, -7, 2, 16, -10, -16, 10, 15, -11, 3, 8, -21, -11, 15, -17, -21, -22, 10, 4, -14, -8, -1, -3, -15, 14, -6, 19, 17, 21, -15, 13, -15, -18, 17, 2, -3, -19, -47, -44, -33, -60, -45, -20, -22, -32, 6, 21, -1, 6, 17, 6, 14, 14, 1, 19, 9, -20, 8, -18, 17, -4, -19, 44, -77, -77, -53, -44, -83, -81, -58, -77, -68, -33, -40, 44, 24, 24, 19, 3, 5, -13, -9, 5, -14, -4, -20, 0, 16, 10, 47, -5, -95, -85, -77, -96, -89, -81, -91, -85, -97, -67, -26, -20, 16, 11, -13, -12, -6, 14, -11, -8, 15, -7, 7, 25, -6, 21, 41, 32, -39, -61, -40, -43, -73, -89, -129, -112, -94, -95, -37, -27, 4, -4, 5, 7, 20, -11, -9, 17, -12, -19, -1, 19, 51, 24, 34, 5, -84, -58, -52, -50, -102, -89, -115, -85, -95, -69, -21, 12, 8, 18, 3, -20, 12, 4, 19, -17, 17, -20, 40, 47, 49, 27, 5, -7, -18, -37, -27, -47, -80, -63, -97, -71, -46, -17, 32, 39, -26, -41, 17, 10, -4, -8, -7, 8, 17, 1, 53, 37, 32, -10, -15, -1, 4, 8, 13, -11, -10, -30, -60, -35, -27, -15, 33, 68, 72, 14, 6, 15, 11, -6, 0, 19, 10, -14, 18, -18, 31, 1, 17, 19, -16, -32, -13, 2, -10, -14, -33, -32, -13, -17, 11, 62, 67, -21, -37, -25, -9, 16, -6, 16, 1, 19, 20, -58, 9, 12, -3, 7, 5, 17, 4, -1, 24, -3, -28, 5, -20, -9, 9, 61, 54, -13, -3, 14, -4, 6, 10, 10, 6, -8, -8, -18, -10, -5, -6, 0, 22, 12, -5, -17, -3, 6, 6, 26, 8, 13, 53, 73, 63, -17, 26, 57, 7, 10, 17, -4, -16, 8, -29, -4, 16, -43, -42, -37, -20, -40, -24, -9, -31, 20, 32, 46, 41, 38, 79, 84, 22, 34, 2, 22, 1, -17, -18, -16, -9, 1, -2, 47, 21, -18, -50, -47, -21, -35, -13, 11, 32, 57, 42, 53, 70, 82, 76, 64, 25, 14, -11, 65, 9, -12, 14, -3, 18, 12, 44, 65, 9, 5, 10, 17, 15, 1, 25, 40, 30, 71, 51, 58, 53, 69, 27, 28, -8, -12, -16, 33, -10, 15, -4, -2, 27, 0, 27, 52, 28, 13, 27, -2, 11, -16, 17, 19, 4, 19, 41, 28, 38, 13, 17, -24, -27, -50, -11, 26, 6, -2, 7, 19, -4, -1, 11, 27, 4, 9, 3, -3, 4, 15, 27, 31, 38, 44, 44, 33, 19, -3, -7, -40, -62, -61, -44, 11, 9, 4, 18, -17, 32, -11, 13, 30, 39, 15, 42, 23, 36, 31, 53, 41, 34, -3, -1, 24, 2, -21, -10, -31, -66, -38, -56, 18, 14, 5, 5, 8, 0, -8, -19, 37, 29, 13, 47, 0, 11, -3, 20, 35, 26, -32, -5, -9, -35, -17, -11, -22, -35, -1, -31, 9, 20, 11, -3, 20, -13, 2, -8, 26, 4, 16, -12, -51, -59, -50, 12, 37, -8, -18, -17, -9, -10, -50, -30, -14, -33, -36, -59, 51, 19, 21, -13, -15, 17, -30, -21, -8, -49, -63, -55, -2, -39, -2, -10, -5, -17, -10, -11, -2, -14, -37, -25, -21, -32, 23, -35, 37, -18, 8, 18, 19, 3, -24, -3, 0, -13, -28, -42, -51, -13, 20, 42, 18, 15, -7, -36, -34, -7, -37, -40, -58, -49, -40, -10, 20, -3, -7, 14, 0, -7, -37, 1, -10, -10, -29, 1, 4, -33, -4, 5, -6, -20, -25, -38, -14, 10, -38, -44, -13, -8, -25, -19, 19, -1, 12, 14, 13, 16, -2, -8, -28, -47, -60, -55, -43, 9, -3, 21, 23, -11, -20, -21, -27, -27, -39, -29, -47, 0, -17, -34, -3, -18, 0, 2, -13, 13, -1, 40, 0, -22, -40, -72, -39, -14, -1, 21, 13, 2, 11, -14, -51, -38, -33, -38, -13, -2, -24, -19, -22, 20, 14, -4, 10, 7, 17, 24, 31, 31, -18, -22, -32, -1, -6, 21, 36, -35, -9, -52, -30, -36, -9, 2, -21, -20, -36, -22, -13, -19, -7, 3, 11, -19, -21, 43, 17, 0, 9, -14, -14, -23, -4, 31, 27, 41, 17, 32, -3, -14, 13, 2, 10, 8, -41, -26, -38, -9, 14, 1, -1, 2, -32, -5, -29, -6, -14, -7, -7, 17, -37, 29, 6, 1, 31, -10, -2, -18, -24, -25, -44, -32, -57, -42, 2),
  125 => (-17, -7, 1, 9, 3, -2, 15, 10, -2, -5, 9, -15, 10, -4, -19, 15, 3, -16, 34, 12, 1, 7, 9, 4, -14, 14, 4, -3, 18, -19, -18, -1, -8, -14, -2, 14, 3, -9, -6, 1, 1, -4, 24, -22, 38, -9, 10, 12, -17, 10, -12, 6, 14, -3, -8, 15, -6, 17, -8, 1, 4, -7, 17, -18, -10, 12, 9, 39, -5, -19, -17, 0, -41, -48, -18, -24, -25, 4, -16, 10, -12, -13, -15, 18, -15, -18, -12, -18, 0, 20, 3, -16, 11, 45, -6, 4, 53, 56, 45, 33, -72, -65, -68, -42, -16, -4, -10, -28, -11, 16, -13, 13, -13, -2, -17, 13, -12, 20, -14, -10, 5, -24, -28, -8, 56, 66, 50, -14, -66, -67, -70, -26, -61, -20, -35, -21, 1, 15, 15, -7, -7, 5, -4, -9, 3, -6, 11, -21, -14, -82, -81, 10, 64, 73, -4, -19, -56, -67, -29, -25, -18, 7, 0, 14, -7, -6, 3, 15, 4, -18, 20, -3, -15, -5, -13, -10, -46, -143, -63, 16, 44, -12, -12, -31, -63, -15, -10, -5, 8, 35, 34, 26, 12, -24, 14, 1, 18, -19, 5, -2, 5, -19, -15, -25, -65, -137, -58, 39, 1, -20, 1, -22, -16, 2, 11, 24, 43, 25, 27, 11, -14, 3, 1, -18, -19, -16, -14, -10, 19, 1, -23, -32, -48, -97, -21, 13, -20, -15, -6, -53, -34, 1, -31, 9, 5, 12, -33, -35, 0, -32, 9, 11, 17, -6, -7, 16, -7, 6, -52, -16, -59, -95, -16, 17, 15, -16, -20, -40, -35, -1, 16, -14, 1, -32, -19, -75, -25, -24, -7, -11, -7, 15, -14, -14, -2, -3, -22, -49, -48, -61, -16, -13, -10, -17, -39, -38, -38, -36, -40, -31, -36, -49, -70, -73, -27, -40, 1, 18, 21, 10, 17, 15, 20, 11, -28, -40, -39, 17, 20, 9, -5, -21, -76, -87, -104, -93, -71, -67, -53, -20, -72, -148, -41, -7, -35, 15, 6, -5, 12, -11, 0, -20, -16, -22, 1, 35, 72, 23, 30, 33, -21, -18, -21, -56, -67, -60, -60, -45, -99, -89, -81, -43, -23, 1, 19, -7, 9, -3, -6, 17, 8, 6, 31, 71, 69, 45, 53, 21, 17, 8, 40, -3, 0, 7, 16, -6, -50, -70, -41, -14, 35, 49, 4, 18, -8, -11, 6, -7, 12, 14, -13, 30, 28, 18, 28, 22, 8, 15, 0, -16, 23, 17, -3, 16, 3, -21, -7, 19, 11, 56, -6, 14, -15, 5, -36, 2, 36, -8, -18, 10, 7, -4, 29, 13, -3, 28, 9, -2, 8, 29, 13, 24, 13, 43, -1, 20, 8, 26, 10, -2, 7, 9, -1, 0, 24, 59, 10, -6, -26, 14, 15, -17, 4, 24, 9, -4, -14, 19, 27, 33, 32, 29, 44, 15, 31, -1, 12, 8, -17, -18, -7, 31, 24, 39, 26, -4, 2, 3, 10, 7, -9, -1, 8, -7, 13, 12, 30, 28, 32, 40, 51, 28, 52, 19, 17, -6, -9, -6, 0, -27, 9, -14, 6, -9, 9, 20, 33, -10, -21, 6, -16, -3, 8, 32, 35, 48, 42, 28, 63, 31, 7, -9, -13, 14, -3, 20, 13, -24, -29, -46, -13, -12, 19, 29, 10, 7, 0, -13, -40, -19, -6, 13, 41, 40, 35, 79, 71, 32, -8, 12, 3, -4, -10, 0, -21, -45, -21, -37, -5, 30, 31, 33, 26, 16, 0, -2, -13, -12, 23, 32, 17, 22, 52, 46, 59, 33, 32, 6, 18, 0, 18, -1, -12, -40, -39, -33, 6, 12, 14, 23, 4, 40, 20, -13, 11, -10, 29, 35, 3, -8, 16, 14, 40, 46, 6, 6, -4, -18, 14, 11, -11, -84, -49, -41, -16, 12, 30, -2, 23, 16, 8, -5, 6, 25, -2, -1, 12, -12, -2, 8, 15, 38, 11, -31, 13, 18, 15, 11, -10, -48, -47, -54, -35, -50, -1, -3, -31, 1, 10, 31, -13, -5, 11, -11, -33, 2, 22, 27, 29, 37, 26, -2, 12, 3, 16, -6, 1, -24, -52, -57, -48, -28, -43, -34, -55, -22, -2, -20, 2, -34, -21, -34, -24, -33, -3, 20, 10, 3, 14, 9, -5, -11, -3, 1, -18, -1, -15, -32, 3, -52, -35, 0, -48, -31, -28, -37, -76, -55, -51, -30, -17, -34, -10, -12, 7, 12, -17, 33, 13, -20, -5, -4, 8, -5, 7, -20, -7, -6, -25, 15, -20, -23, -22, -52, -58, -41, -28, -41, -52, -42, -18, -10, -13, 13, -26, 11, -8, 16, 12, 17, 5, -20, 3, -6, -25, -21, 3, 4, -7, 25, -18, -31, -44, -58, -51, -48, -75, -17, -40, 1, -17, 2, -35, 11),
  126 => (-17, -1, 4, -5, -18, -12, -14, -10, -15, 1, -19, -8, -10, -19, -23, 8, -40, -34, -38, -75, -96, -39, -28, 16, -19, -13, -17, 14, -2, -8, -8, 9, -9, 0, 11, 14, 21, 19, -6, 13, 16, -8, 34, 49, 49, 45, 27, 48, 46, 25, 31, -28, -5, -2, 9, 9, 1, 14, 10, 6, 4, 14, 13, -11, -17, -12, -25, -1, 30, 21, 10, -16, -4, 11, 30, 16, 55, 62, 40, 9, 4, -11, -11, -19, -16, -2, -2, 7, -18, 6, 17, -2, 21, -29, -32, -1, 22, -27, 7, -3, -24, -5, 18, 19, 17, 52, 67, 48, -3, 31, -17, 13, -3, -10, -2, -4, 3, -10, 4, -2, 1, -43, -9, 33, -4, 10, -2, 4, -9, 6, 8, 4, -1, 40, 29, -1, -31, -10, -12, -1, -4, -20, 4, 15, -3, -1, -29, 13, -12, -16, 25, 24, 28, 8, -9, -27, -15, 10, 18, 12, -7, -4, -40, -15, -41, -2, -7, 4, 11, -10, 8, -12, 4, 1, -42, -14, -34, 22, 37, 7, 22, 28, -9, -27, -29, 20, -9, -21, -4, -27, -31, -41, -53, 11, -8, -19, -14, -15, 8, 13, -3, 11, 3, 18, 67, 58, 12, 5, 10, 48, -7, -2, 11, -13, -3, -17, 45, 16, -16, -50, -51, -39, 14, 31, 4, 15, -20, -2, -2, -19, 8, 57, 55, 69, 37, 2, 47, -4, -5, 16, 2, 5, 30, -29, -3, 8, -38, 2, 18, 46, 23, 37, 19, -1, 6, -17, -10, 2, 7, 59, 95, 78, 56, 63, 31, 51, 29, 41, -2, 11, 21, 12, 32, 15, 14, -11, 48, 61, 59, 89, 6, -18, -8, -2, 19, 10, 49, 83, 91, 90, 76, 74, 71, 36, 70, 60, 53, 48, 37, -1, 62, 37, -14, 23, 27, 41, 59, 23, -7, 15, 18, -13, 20, 0, 39, 57, 69, 102, 89, 48, 55, 37, 83, 97, 78, 68, 42, 55, 58, 16, 11, 6, 16, 18, 77, 29, -6, -17, 8, -16, 18, 3, 48, 65, 52, 75, 73, 11, 29, 20, 65, 83, 53, 64, 39, 22, 28, 23, 11, -2, 23, 52, 67, 27, 17, 10, -9, -2, -25, -7, 35, 55, 42, 41, 50, 61, 54, 22, 49, 27, 55, 52, 32, 21, 40, 28, 45, 7, 40, 12, 84, 50, -5, -18, 14, 12, -38, 13, 17, -1, 20, 18, 19, 33, 35, 42, 45, 50, 48, 52, 49, 66, 48, 46, 12, -6, 57, 34, 65, 44, -2, 1, 0, 3, -19, 24, 41, 13, -3, -17, 33, 53, 6, 4, 4, 43, 42, 32, 56, 45, 60, 30, -4, -12, 22, 42, 18, 0, -16, -19, 20, 3, 24, 26, 44, -6, -25, -12, 10, 6, -3, 16, -7, 32, 15, 8, 53, 50, 39, -5, 11, -8, 12, 3, 5, 2, 9, 5, 4, 19, 41, -12, -23, -54, 6, 4, -24, -28, -2, 10, 47, 31, 21, 20, 6, 13, 1, 5, 30, 19, 0, 14, 19, 47, 12, -2, -18, -14, 4, -19, -43, -56, -13, -42, -57, -13, 15, 17, 53, 8, 10, 20, 28, 7, 6, 8, 27, 33, 11, 20, 52, 10, -4, -3, -10, -15, -15, 25, -9, -38, -43, -27, -80, -36, -1, 21, -7, 12, 21, -3, 19, 10, 25, 8, 6, 34, 29, 1, 17, -20, -2, 11, 20, -3, 30, 30, 9, -41, -47, -47, -55, -43, 0, -6, -17, 5, 16, 1, -13, -1, 23, 6, 28, 22, 23, 31, 34, -11, -7, 15, 15, -18, 6, 29, 4, -33, 1, -17, 15, -1, -37, -26, -29, 0, -3, -10, 3, -5, -26, -28, -15, -3, 58, 3, 24, -15, 13, -8, -2, 0, -16, 32, -4, 4, -40, -57, -30, -15, -14, -31, -24, 1, 4, 30, 22, -3, -19, -15, -25, 13, 32, -29, -33, -35, -13, -16, 6, 13, -15, 10, -6, 16, -21, -28, 11, 20, -15, 11, 6, 32, 19, 42, 35, -2, -19, 11, 29, 12, 0, -5, -7, -38, -12, 14, -16, -5, -10, -10, -13, 13, -13, 6, 33, 20, -7, 13, 21, 8, -2, 23, 8, -20, -18, -6, 9, 39, 30, 22, 2, -29, -19, 14, -15, -15, 23, -6, -2, -9, 10, -37, 17, -4, -24, -12, 16, 19, -16, 16, 5, -6, -11, -21, -26, 1, 47, 60, 19, -44, -10, -8, -8, -15, -24, 8, 8, -5, 5, 19, 47, 1, 16, 27, -2, 28, -3, 14, -17, -42, -20, -8, -3, -31, 31, 44, -25, -23, 12, 21, -1, -13, 20, 28, 58, 52, 72, 42, 61, 64, 62, 42, 64, 58, 54, 61, -12, -9, 7, 16, 20, -19, -1, 38, -34, -42),
  127 => (-20, -20, -16, -6, 6, 16, -17, -8, -2, 17, 16, -5, 15, 3, 24, 18, 29, 10, 0, 5, 11, -17, -30, 2, 2, 20, 17, -8, -6, 18, 5, -6, -18, 10, -5, -11, 5, -12, 21, 0, -39, 8, -28, -16, -30, -6, -26, -22, -10, -50, -16, -25, -35, 3, 7, -2, 20, -6, -4, -5, 14, -4, 4, -8, -4, 2, 5, -25, -42, -15, 40, 72, 67, 57, 45, 1, -32, -40, -70, -41, -28, -11, -14, -13, -14, -20, 8, -7, -9, 11, 2, -9, -13, -25, -21, -12, -5, 34, 54, 67, 36, 70, 43, 50, -10, -25, -16, -11, -41, 24, -18, 19, -10, -14, 17, -16, -7, 16, 9, -15, -53, -29, -45, 4, -8, 51, 55, 48, 65, 36, 6, -13, 0, -37, -31, -20, -33, -33, 17, 11, 6, -15, -17, -19, 14, -5, -25, -44, -67, -80, -44, -15, 14, -3, 35, 26, 4, -8, -25, -41, -23, 4, -26, 11, -21, -18, -9, -18, 11, 14, -9, -18, 5, -1, -50, -63, -67, -33, -14, 13, 6, 17, 14, 34, -14, 26, 10, 2, 2, 28, 12, 35, 1, 2, 5, 0, -9, 12, -18, 20, 15, -6, -45, -76, -73, -11, 33, -25, -19, -7, -5, 59, 2, 3, 14, 13, 59, 24, 2, 52, 47, -9, 75, 12, -18, 11, -1, -19, 19, 8, -54, -28, -23, -17, -25, -53, -76, -43, -8, 29, 32, 18, 29, 42, 19, 33, -8, 24, 35, 56, 61, 37, -5, -11, 3, 0, 8, -9, 1, 20, -30, -19, -45, -47, -45, -52, 3, 40, 54, 45, 63, 37, 65, 38, -8, 9, 32, 38, 24, 87, -17, -3, 18, 1, -19, 25, 22, 42, 6, 14, -10, 1, 25, 3, -15, 44, 56, 46, 66, 77, 84, 48, 14, 7, 5, 53, 62, 59, 6, 7, 6, 8, -1, 42, 113, 40, 70, 59, 49, 39, 61, 62, 36, 58, 50, 47, 25, 39, 51, 32, 32, 39, 32, 38, 55, 73, 5, -9, -10, -19, -12, 62, 125, 81, 63, 66, 84, 73, 61, 62, 40, 78, 43, 46, 23, 52, 10, 17, 37, 23, 13, 78, 48, 44, 14, -18, 15, 20, -7, 31, 76, 75, 72, 56, 50, 50, 31, 8, 34, 23, 28, 36, 17, 15, 59, 23, 39, 46, 39, 35, 33, 10, 17, -9, -4, 4, -14, 53, 69, 44, 52, 25, 17, 20, 6, 2, 8, 1, 72, 58, 22, 13, 20, -9, 12, 34, 37, 61, 37, -3, 20, 5, 20, -10, 13, 18, 40, 36, 61, 53, 42, 35, 45, 38, 11, 32, 22, 14, 7, 18, 27, -29, -11, 5, -1, 40, -20, -17, -17, 20, 18, 8, 39, 20, 65, 41, 45, 36, 8, 23, 53, 37, 33, 32, 13, -6, -10, 19, 35, 0, 27, -6, -46, -16, -12, -45, -8, 15, -15, -6, 28, 19, 45, 27, 46, 29, 29, 11, 10, 46, 14, 17, 2, -5, -7, 4, 32, 12, 3, 18, -14, 34, 19, -3, -7, -3, -17, -7, 5, 2, 23, 1, -5, 24, 21, 2, 6, 11, 30, 17, 23, -16, -30, -41, -5, -16, -21, 1, -12, 5, 19, -1, 11, 8, 12, 10, 13, -19, 24, -26, 30, 30, 8, 1, 43, 0, -12, 4, 3, 9, -22, -2, -47, -4, -18, 7, -14, 15, 11, 38, 13, -12, 8, 8, -43, -45, -21, -7, 16, 13, -2, -25, 3, -5, -24, -52, -20, -27, 17, 10, 11, -19, -25, -27, -3, 13, 11, -35, -17, 20, -6, -20, -36, -37, -11, 3, -14, -7, -21, -48, -27, -13, -30, -19, -6, 12, -6, 5, -14, -25, -1, 7, -1, 15, -9, -3, -13, 1, 11, 7, -23, -18, -15, 15, 11, -19, -36, -44, -50, -33, -43, -14, -15, 15, 12, 25, 27, -36, -29, -16, -2, 8, -31, -58, 8, 5, 10, 21, -23, -32, -52, 7, -15, -23, -35, -19, -24, -7, -60, -27, -18, 18, 20, 13, 6, -25, -37, -14, 3, 13, -14, -37, -9, 12, -9, 13, -37, -31, -32, -9, 8, -33, -26, -38, -29, -18, -37, -44, -17, -14, 1, -2, 5, 12, -29, 29, 17, 57, 25, -8, 16, -10, 12, 10, -18, -27, -20, -30, -13, -8, 27, 17, -7, 19, 8, -10, -17, 25, 24, 18, 2, 8, -5, 53, 16, 19, 17, -23, 19, -3, 12, 6, -13, -32, -46, -28, 1, 23, 55, -10, -3, 23, 29, 27, 22, 20, 28, -9, -3, -7, -2, 20, -16, 0, 5, -44, -2, -18, -2, -8, -15, -25, -28, -47, -26, -39, -29, -35, -2, 5, 3, -33, -10, 18, -17, -47, -41, -69, -55, -53, -27, -28, -57, -12)
);
end package;

package body Layer1_Weights is
end package body;