library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.Types.all;


entity Top_tb is
end Top_tb;

architecture behavior of Top_tb is

    -- Bileşeni test edilecek üst modül
    component Top
        Port (
            clk    : in  std_logic;
			input_data : in  integer_vector(0 to 783);
            result : out integer;
			layer6_out  : out integer_vector(0 to 9);
			layer1_out_dbg  : out integer_vector(0 to 127);
			layer4_out_dbg  : out integer_vector(0 to 63)
        );
    end component;

    -- Testbench sinyalleri
    signal clk_tb     : std_logic := '0';
	signal input_data_tb : integer_vector(0 to 783) := (others => 0);
	signal layer1_out_dbg : integer_vector(0 to 127);
	signal layer4_out_dbg : integer_vector(0 to 63);
	signal layer6_out : integer_vector(0 to 9);
    signal result_tb  : integer;

begin

    -- DUT (Device Under Test) instance
    uut: Top
        port map (
            clk    => clk_tb,
			input_data => input_data_tb,
            result => result_tb,
			layer1_out_dbg => layer1_out_dbg,
			layer4_out_dbg => layer4_out_dbg,
			layer6_out  => layer6_out
        );

    -- Saat üretimi: 10 ns periyot
    clk_process : process
    begin
        while now < 2000 ns loop
            clk_tb <= '0';
            wait for 5 ns;
            clk_tb <= '1';
            wait for 5 ns;
        end loop;
        wait;
    end process;
	
    stimulus : process
    begin
        wait for 10 ns;
			input_data_tb(0) <= 0;
			input_data_tb(1) <= 0;
			input_data_tb(2) <= 0;
			input_data_tb(3) <= 0;
			input_data_tb(4) <= 0;
			input_data_tb(5) <= 0;
			input_data_tb(6) <= 0;
			input_data_tb(7) <= 0;
			input_data_tb(8) <= 0;
			input_data_tb(9) <= 0;
			input_data_tb(10) <= 0;
			input_data_tb(11) <= 0;
			input_data_tb(12) <= 0;
			input_data_tb(13) <= 0;
			input_data_tb(14) <= 0;
			input_data_tb(15) <= 0;
			input_data_tb(16) <= 0;
			input_data_tb(17) <= 0;
			input_data_tb(18) <= 0;
			input_data_tb(19) <= 0;
			input_data_tb(20) <= 0;
			input_data_tb(21) <= 0;
			input_data_tb(22) <= 0;
			input_data_tb(23) <= 0;
			input_data_tb(24) <= 0;
			input_data_tb(25) <= 0;
			input_data_tb(26) <= 0;
			input_data_tb(27) <= 0;
			input_data_tb(28) <= 0;
			input_data_tb(29) <= 0;
			input_data_tb(30) <= 0;
			input_data_tb(31) <= 0;
			input_data_tb(32) <= 0;
			input_data_tb(33) <= 0;
			input_data_tb(34) <= 0;
			input_data_tb(35) <= 0;
			input_data_tb(36) <= 0;
			input_data_tb(37) <= 0;
			input_data_tb(38) <= 0;
			input_data_tb(39) <= 0;
			input_data_tb(40) <= 0;
			input_data_tb(41) <= 0;
			input_data_tb(42) <= 0;
			input_data_tb(43) <= 0;
			input_data_tb(44) <= 0;
			input_data_tb(45) <= 0;
			input_data_tb(46) <= 0;
			input_data_tb(47) <= 0;
			input_data_tb(48) <= 0;
			input_data_tb(49) <= 0;
			input_data_tb(50) <= 0;
			input_data_tb(51) <= 0;
			input_data_tb(52) <= 0;
			input_data_tb(53) <= 0;
			input_data_tb(54) <= 0;
			input_data_tb(55) <= 0;
			input_data_tb(56) <= 0;
			input_data_tb(57) <= 0;
			input_data_tb(58) <= 0;
			input_data_tb(59) <= 0;
			input_data_tb(60) <= 0;
			input_data_tb(61) <= 0;
			input_data_tb(62) <= 0;
			input_data_tb(63) <= 0;
			input_data_tb(64) <= 0;
			input_data_tb(65) <= 0;
			input_data_tb(66) <= 0;
			input_data_tb(67) <= 0;
			input_data_tb(68) <= 0;
			input_data_tb(69) <= 0;
			input_data_tb(70) <= 0;
			input_data_tb(71) <= 0;
			input_data_tb(72) <= 0;
			input_data_tb(73) <= 0;
			input_data_tb(74) <= 0;
			input_data_tb(75) <= 0;
			input_data_tb(76) <= 0;
			input_data_tb(77) <= 0;
			input_data_tb(78) <= 0;
			input_data_tb(79) <= 0;
			input_data_tb(80) <= 0;
			input_data_tb(81) <= 0;
			input_data_tb(82) <= 0;
			input_data_tb(83) <= 0;
			input_data_tb(84) <= 0;
			input_data_tb(85) <= 0;
			input_data_tb(86) <= 0;
			input_data_tb(87) <= 0;
			input_data_tb(88) <= 0;
			input_data_tb(89) <= 0;
			input_data_tb(90) <= 0;
			input_data_tb(91) <= 0;
			input_data_tb(92) <= 0;
			input_data_tb(93) <= 0;
			input_data_tb(94) <= 0;
			input_data_tb(95) <= 0;
			input_data_tb(96) <= 0;
			input_data_tb(97) <= 0;
			input_data_tb(98) <= 0;
			input_data_tb(99) <= 0;
			input_data_tb(100) <= 0;
			input_data_tb(101) <= 0;
			input_data_tb(102) <= 0;
			input_data_tb(103) <= 0;
			input_data_tb(104) <= 0;
			input_data_tb(105) <= 0;
			input_data_tb(106) <= 0;
			input_data_tb(107) <= 0;
			input_data_tb(108) <= 0;
			input_data_tb(109) <= 0;
			input_data_tb(110) <= 0;
			input_data_tb(111) <= 0;
			input_data_tb(112) <= 0;
			input_data_tb(113) <= 0;
			input_data_tb(114) <= 0;
			input_data_tb(115) <= 0;
			input_data_tb(116) <= 0;
			input_data_tb(117) <= 0;
			input_data_tb(118) <= 0;
			input_data_tb(119) <= 0;
			input_data_tb(120) <= 0;
			input_data_tb(121) <= 0;
			input_data_tb(122) <= 0;
			input_data_tb(123) <= 0;
			input_data_tb(124) <= 0;
			input_data_tb(125) <= 0;
			input_data_tb(126) <= 0;
			input_data_tb(127) <= 0;
			input_data_tb(128) <= 0;
			input_data_tb(129) <= 0;
			input_data_tb(130) <= 0;
			input_data_tb(131) <= 0;
			input_data_tb(132) <= 0;
			input_data_tb(133) <= 0;
			input_data_tb(134) <= 0;
			input_data_tb(135) <= 0;
			input_data_tb(136) <= 0;
			input_data_tb(137) <= 0;
			input_data_tb(138) <= 0;
			input_data_tb(139) <= 0;
			input_data_tb(140) <= 0;
			input_data_tb(141) <= 0;
			input_data_tb(142) <= 0;
			input_data_tb(143) <= 0;
			input_data_tb(144) <= 0;
			input_data_tb(145) <= 0;
			input_data_tb(146) <= 0;
			input_data_tb(147) <= 0;
			input_data_tb(148) <= 0;
			input_data_tb(149) <= 0;
			input_data_tb(150) <= 0;
			input_data_tb(151) <= 0;
			input_data_tb(152) <= 255;
			input_data_tb(153) <= 255;
			input_data_tb(154) <= 255;
			input_data_tb(155) <= 255;
			input_data_tb(156) <= 255;
			input_data_tb(157) <= 255;
			input_data_tb(158) <= 0;
			input_data_tb(159) <= 0;
			input_data_tb(160) <= 0;
			input_data_tb(161) <= 0;
			input_data_tb(162) <= 0;
			input_data_tb(163) <= 0;
			input_data_tb(164) <= 0;
			input_data_tb(165) <= 0;
			input_data_tb(166) <= 0;
			input_data_tb(167) <= 0;
			input_data_tb(168) <= 0;
			input_data_tb(169) <= 0;
			input_data_tb(170) <= 0;
			input_data_tb(171) <= 0;
			input_data_tb(172) <= 0;
			input_data_tb(173) <= 0;
			input_data_tb(174) <= 0;
			input_data_tb(175) <= 0;
			input_data_tb(176) <= 0;
			input_data_tb(177) <= 0;
			input_data_tb(178) <= 255;
			input_data_tb(179) <= 255;
			input_data_tb(180) <= 255;
			input_data_tb(181) <= 255;
			input_data_tb(182) <= 255;
			input_data_tb(183) <= 255;
			input_data_tb(184) <= 255;
			input_data_tb(185) <= 255;
			input_data_tb(186) <= 255;
			input_data_tb(187) <= 0;
			input_data_tb(188) <= 0;
			input_data_tb(189) <= 0;
			input_data_tb(190) <= 0;
			input_data_tb(191) <= 0;
			input_data_tb(192) <= 0;
			input_data_tb(193) <= 0;
			input_data_tb(194) <= 0;
			input_data_tb(195) <= 0;
			input_data_tb(196) <= 0;
			input_data_tb(197) <= 0;
			input_data_tb(198) <= 0;
			input_data_tb(199) <= 0;
			input_data_tb(200) <= 0;
			input_data_tb(201) <= 0;
			input_data_tb(202) <= 0;
			input_data_tb(203) <= 0;
			input_data_tb(204) <= 0;
			input_data_tb(205) <= 255;
			input_data_tb(206) <= 255;
			input_data_tb(207) <= 255;
			input_data_tb(208) <= 255;
			input_data_tb(209) <= 255;
			input_data_tb(210) <= 255;
			input_data_tb(211) <= 255;
			input_data_tb(212) <= 255;
			input_data_tb(213) <= 255;
			input_data_tb(214) <= 255;
			input_data_tb(215) <= 0;
			input_data_tb(216) <= 0;
			input_data_tb(217) <= 0;
			input_data_tb(218) <= 0;
			input_data_tb(219) <= 0;
			input_data_tb(220) <= 0;
			input_data_tb(221) <= 0;
			input_data_tb(222) <= 0;
			input_data_tb(223) <= 0;
			input_data_tb(224) <= 0;
			input_data_tb(225) <= 0;
			input_data_tb(226) <= 0;
			input_data_tb(227) <= 0;
			input_data_tb(228) <= 0;
			input_data_tb(229) <= 0;
			input_data_tb(230) <= 0;
			input_data_tb(231) <= 0;
			input_data_tb(232) <= 255;
			input_data_tb(233) <= 255;
			input_data_tb(234) <= 255;
			input_data_tb(235) <= 255;
			input_data_tb(236) <= 0;
			input_data_tb(237) <= 0;
			input_data_tb(238) <= 0;
			input_data_tb(239) <= 0;
			input_data_tb(240) <= 255;
			input_data_tb(241) <= 255;
			input_data_tb(242) <= 255;
			input_data_tb(243) <= 255;
			input_data_tb(244) <= 0;
			input_data_tb(245) <= 0;
			input_data_tb(246) <= 0;
			input_data_tb(247) <= 0;
			input_data_tb(248) <= 0;
			input_data_tb(249) <= 0;
			input_data_tb(250) <= 0;
			input_data_tb(251) <= 0;
			input_data_tb(252) <= 0;
			input_data_tb(253) <= 0;
			input_data_tb(254) <= 0;
			input_data_tb(255) <= 0;
			input_data_tb(256) <= 0;
			input_data_tb(257) <= 0;
			input_data_tb(258) <= 0;
			input_data_tb(259) <= 255;
			input_data_tb(260) <= 255;
			input_data_tb(261) <= 255;
			input_data_tb(262) <= 255;
			input_data_tb(263) <= 0;
			input_data_tb(264) <= 0;
			input_data_tb(265) <= 0;
			input_data_tb(266) <= 0;
			input_data_tb(267) <= 0;
			input_data_tb(268) <= 0;
			input_data_tb(269) <= 255;
			input_data_tb(270) <= 255;
			input_data_tb(271) <= 255;
			input_data_tb(272) <= 0;
			input_data_tb(273) <= 0;
			input_data_tb(274) <= 0;
			input_data_tb(275) <= 0;
			input_data_tb(276) <= 0;
			input_data_tb(277) <= 0;
			input_data_tb(278) <= 0;
			input_data_tb(279) <= 0;
			input_data_tb(280) <= 0;
			input_data_tb(281) <= 0;
			input_data_tb(282) <= 0;
			input_data_tb(283) <= 0;
			input_data_tb(284) <= 0;
			input_data_tb(285) <= 0;
			input_data_tb(286) <= 0;
			input_data_tb(287) <= 255;
			input_data_tb(288) <= 255;
			input_data_tb(289) <= 255;
			input_data_tb(290) <= 255;
			input_data_tb(291) <= 0;
			input_data_tb(292) <= 0;
			input_data_tb(293) <= 0;
			input_data_tb(294) <= 0;
			input_data_tb(295) <= 0;
			input_data_tb(296) <= 0;
			input_data_tb(297) <= 255;
			input_data_tb(298) <= 255;
			input_data_tb(299) <= 255;
			input_data_tb(300) <= 0;
			input_data_tb(301) <= 0;
			input_data_tb(302) <= 0;
			input_data_tb(303) <= 0;
			input_data_tb(304) <= 0;
			input_data_tb(305) <= 0;
			input_data_tb(306) <= 0;
			input_data_tb(307) <= 0;
			input_data_tb(308) <= 0;
			input_data_tb(309) <= 0;
			input_data_tb(310) <= 0;
			input_data_tb(311) <= 0;
			input_data_tb(312) <= 0;
			input_data_tb(313) <= 0;
			input_data_tb(314) <= 0;
			input_data_tb(315) <= 0;
			input_data_tb(316) <= 0;
			input_data_tb(317) <= 0;
			input_data_tb(318) <= 0;
			input_data_tb(319) <= 0;
			input_data_tb(320) <= 0;
			input_data_tb(321) <= 0;
			input_data_tb(322) <= 0;
			input_data_tb(323) <= 0;
			input_data_tb(324) <= 0;
			input_data_tb(325) <= 255;
			input_data_tb(326) <= 255;
			input_data_tb(327) <= 255;
			input_data_tb(328) <= 0;
			input_data_tb(329) <= 0;
			input_data_tb(330) <= 0;
			input_data_tb(331) <= 0;
			input_data_tb(332) <= 0;
			input_data_tb(333) <= 0;
			input_data_tb(334) <= 0;
			input_data_tb(335) <= 0;
			input_data_tb(336) <= 0;
			input_data_tb(337) <= 0;
			input_data_tb(338) <= 0;
			input_data_tb(339) <= 0;
			input_data_tb(340) <= 0;
			input_data_tb(341) <= 0;
			input_data_tb(342) <= 0;
			input_data_tb(343) <= 0;
			input_data_tb(344) <= 0;
			input_data_tb(345) <= 0;
			input_data_tb(346) <= 0;
			input_data_tb(347) <= 0;
			input_data_tb(348) <= 0;
			input_data_tb(349) <= 0;
			input_data_tb(350) <= 0;
			input_data_tb(351) <= 0;
			input_data_tb(352) <= 0;
			input_data_tb(353) <= 255;
			input_data_tb(354) <= 255;
			input_data_tb(355) <= 255;
			input_data_tb(356) <= 0;
			input_data_tb(357) <= 0;
			input_data_tb(358) <= 0;
			input_data_tb(359) <= 0;
			input_data_tb(360) <= 0;
			input_data_tb(361) <= 0;
			input_data_tb(362) <= 0;
			input_data_tb(363) <= 0;
			input_data_tb(364) <= 0;
			input_data_tb(365) <= 0;
			input_data_tb(366) <= 0;
			input_data_tb(367) <= 0;
			input_data_tb(368) <= 0;
			input_data_tb(369) <= 0;
			input_data_tb(370) <= 0;
			input_data_tb(371) <= 0;
			input_data_tb(372) <= 0;
			input_data_tb(373) <= 0;
			input_data_tb(374) <= 0;
			input_data_tb(375) <= 0;
			input_data_tb(376) <= 0;
			input_data_tb(377) <= 0;
			input_data_tb(378) <= 0;
			input_data_tb(379) <= 0;
			input_data_tb(380) <= 0;
			input_data_tb(381) <= 255;
			input_data_tb(382) <= 255;
			input_data_tb(383) <= 0;
			input_data_tb(384) <= 0;
			input_data_tb(385) <= 0;
			input_data_tb(386) <= 0;
			input_data_tb(387) <= 0;
			input_data_tb(388) <= 0;
			input_data_tb(389) <= 0;
			input_data_tb(390) <= 0;
			input_data_tb(391) <= 0;
			input_data_tb(392) <= 0;
			input_data_tb(393) <= 0;
			input_data_tb(394) <= 0;
			input_data_tb(395) <= 0;
			input_data_tb(396) <= 0;
			input_data_tb(397) <= 0;
			input_data_tb(398) <= 0;
			input_data_tb(399) <= 0;
			input_data_tb(400) <= 0;
			input_data_tb(401) <= 0;
			input_data_tb(402) <= 0;
			input_data_tb(403) <= 0;
			input_data_tb(404) <= 0;
			input_data_tb(405) <= 0;
			input_data_tb(406) <= 0;
			input_data_tb(407) <= 0;
			input_data_tb(408) <= 0;
			input_data_tb(409) <= 255;
			input_data_tb(410) <= 255;
			input_data_tb(411) <= 0;
			input_data_tb(412) <= 0;
			input_data_tb(413) <= 0;
			input_data_tb(414) <= 0;
			input_data_tb(415) <= 0;
			input_data_tb(416) <= 0;
			input_data_tb(417) <= 0;
			input_data_tb(418) <= 0;
			input_data_tb(419) <= 0;
			input_data_tb(420) <= 0;
			input_data_tb(421) <= 0;
			input_data_tb(422) <= 0;
			input_data_tb(423) <= 0;
			input_data_tb(424) <= 0;
			input_data_tb(425) <= 0;
			input_data_tb(426) <= 0;
			input_data_tb(427) <= 0;
			input_data_tb(428) <= 0;
			input_data_tb(429) <= 0;
			input_data_tb(430) <= 0;
			input_data_tb(431) <= 0;
			input_data_tb(432) <= 0;
			input_data_tb(433) <= 0;
			input_data_tb(434) <= 0;
			input_data_tb(435) <= 0;
			input_data_tb(436) <= 255;
			input_data_tb(437) <= 255;
			input_data_tb(438) <= 0;
			input_data_tb(439) <= 0;
			input_data_tb(440) <= 0;
			input_data_tb(441) <= 0;
			input_data_tb(442) <= 0;
			input_data_tb(443) <= 0;
			input_data_tb(444) <= 0;
			input_data_tb(445) <= 0;
			input_data_tb(446) <= 0;
			input_data_tb(447) <= 0;
			input_data_tb(448) <= 0;
			input_data_tb(449) <= 0;
			input_data_tb(450) <= 0;
			input_data_tb(451) <= 0;
			input_data_tb(452) <= 0;
			input_data_tb(453) <= 0;
			input_data_tb(454) <= 0;
			input_data_tb(455) <= 0;
			input_data_tb(456) <= 0;
			input_data_tb(457) <= 0;
			input_data_tb(458) <= 0;
			input_data_tb(459) <= 0;
			input_data_tb(460) <= 0;
			input_data_tb(461) <= 0;
			input_data_tb(462) <= 0;
			input_data_tb(463) <= 255;
			input_data_tb(464) <= 255;
			input_data_tb(465) <= 255;
			input_data_tb(466) <= 0;
			input_data_tb(467) <= 0;
			input_data_tb(468) <= 0;
			input_data_tb(469) <= 0;
			input_data_tb(470) <= 0;
			input_data_tb(471) <= 0;
			input_data_tb(472) <= 0;
			input_data_tb(473) <= 0;
			input_data_tb(474) <= 0;
			input_data_tb(475) <= 0;
			input_data_tb(476) <= 0;
			input_data_tb(477) <= 0;
			input_data_tb(478) <= 0;
			input_data_tb(479) <= 0;
			input_data_tb(480) <= 0;
			input_data_tb(481) <= 0;
			input_data_tb(482) <= 0;
			input_data_tb(483) <= 0;
			input_data_tb(484) <= 0;
			input_data_tb(485) <= 0;
			input_data_tb(486) <= 0;
			input_data_tb(487) <= 0;
			input_data_tb(488) <= 0;
			input_data_tb(489) <= 0;
			input_data_tb(490) <= 255;
			input_data_tb(491) <= 255;
			input_data_tb(492) <= 255;
			input_data_tb(493) <= 0;
			input_data_tb(494) <= 0;
			input_data_tb(495) <= 0;
			input_data_tb(496) <= 0;
			input_data_tb(497) <= 0;
			input_data_tb(498) <= 0;
			input_data_tb(499) <= 0;
			input_data_tb(500) <= 0;
			input_data_tb(501) <= 0;
			input_data_tb(502) <= 0;
			input_data_tb(503) <= 0;
			input_data_tb(504) <= 0;
			input_data_tb(505) <= 0;
			input_data_tb(506) <= 0;
			input_data_tb(507) <= 0;
			input_data_tb(508) <= 0;
			input_data_tb(509) <= 0;
			input_data_tb(510) <= 0;
			input_data_tb(511) <= 0;
			input_data_tb(512) <= 0;
			input_data_tb(513) <= 0;
			input_data_tb(514) <= 0;
			input_data_tb(515) <= 0;
			input_data_tb(516) <= 255;
			input_data_tb(517) <= 255;
			input_data_tb(518) <= 255;
			input_data_tb(519) <= 255;
			input_data_tb(520) <= 0;
			input_data_tb(521) <= 0;
			input_data_tb(522) <= 0;
			input_data_tb(523) <= 0;
			input_data_tb(524) <= 0;
			input_data_tb(525) <= 0;
			input_data_tb(526) <= 0;
			input_data_tb(527) <= 0;
			input_data_tb(528) <= 0;
			input_data_tb(529) <= 0;
			input_data_tb(530) <= 0;
			input_data_tb(531) <= 0;
			input_data_tb(532) <= 0;
			input_data_tb(533) <= 0;
			input_data_tb(534) <= 0;
			input_data_tb(535) <= 0;
			input_data_tb(536) <= 0;
			input_data_tb(537) <= 0;
			input_data_tb(538) <= 0;
			input_data_tb(539) <= 0;
			input_data_tb(540) <= 0;
			input_data_tb(541) <= 0;
			input_data_tb(542) <= 0;
			input_data_tb(543) <= 255;
			input_data_tb(544) <= 255;
			input_data_tb(545) <= 255;
			input_data_tb(546) <= 255;
			input_data_tb(547) <= 0;
			input_data_tb(548) <= 0;
			input_data_tb(549) <= 0;
			input_data_tb(550) <= 0;
			input_data_tb(551) <= 0;
			input_data_tb(552) <= 0;
			input_data_tb(553) <= 0;
			input_data_tb(554) <= 0;
			input_data_tb(555) <= 0;
			input_data_tb(556) <= 0;
			input_data_tb(557) <= 0;
			input_data_tb(558) <= 0;
			input_data_tb(559) <= 0;
			input_data_tb(560) <= 0;
			input_data_tb(561) <= 0;
			input_data_tb(562) <= 0;
			input_data_tb(563) <= 0;
			input_data_tb(564) <= 0;
			input_data_tb(565) <= 0;
			input_data_tb(566) <= 0;
			input_data_tb(567) <= 0;
			input_data_tb(568) <= 255;
			input_data_tb(569) <= 255;
			input_data_tb(570) <= 255;
			input_data_tb(571) <= 255;
			input_data_tb(572) <= 255;
			input_data_tb(573) <= 255;
			input_data_tb(574) <= 255;
			input_data_tb(575) <= 255;
			input_data_tb(576) <= 255;
			input_data_tb(577) <= 255;
			input_data_tb(578) <= 255;
			input_data_tb(579) <= 255;
			input_data_tb(580) <= 255;
			input_data_tb(581) <= 255;
			input_data_tb(582) <= 255;
			input_data_tb(583) <= 255;
			input_data_tb(584) <= 0;
			input_data_tb(585) <= 0;
			input_data_tb(586) <= 0;
			input_data_tb(587) <= 0;
			input_data_tb(588) <= 0;
			input_data_tb(589) <= 0;
			input_data_tb(590) <= 0;
			input_data_tb(591) <= 0;
			input_data_tb(592) <= 255;
			input_data_tb(593) <= 255;
			input_data_tb(594) <= 255;
			input_data_tb(595) <= 255;
			input_data_tb(596) <= 255;
			input_data_tb(597) <= 255;
			input_data_tb(598) <= 255;
			input_data_tb(599) <= 255;
			input_data_tb(600) <= 255;
			input_data_tb(601) <= 255;
			input_data_tb(602) <= 255;
			input_data_tb(603) <= 255;
			input_data_tb(604) <= 255;
			input_data_tb(605) <= 255;
			input_data_tb(606) <= 255;
			input_data_tb(607) <= 255;
			input_data_tb(608) <= 255;
			input_data_tb(609) <= 255;
			input_data_tb(610) <= 255;
			input_data_tb(611) <= 255;
			input_data_tb(612) <= 0;
			input_data_tb(613) <= 0;
			input_data_tb(614) <= 0;
			input_data_tb(615) <= 0;
			input_data_tb(616) <= 0;
			input_data_tb(617) <= 0;
			input_data_tb(618) <= 0;
			input_data_tb(619) <= 0;
			input_data_tb(620) <= 255;
			input_data_tb(621) <= 255;
			input_data_tb(622) <= 255;
			input_data_tb(623) <= 255;
			input_data_tb(624) <= 255;
			input_data_tb(625) <= 255;
			input_data_tb(626) <= 255;
			input_data_tb(627) <= 255;
			input_data_tb(628) <= 255;
			input_data_tb(629) <= 255;
			input_data_tb(630) <= 0;
			input_data_tb(631) <= 255;
			input_data_tb(632) <= 255;
			input_data_tb(633) <= 255;
			input_data_tb(634) <= 255;
			input_data_tb(635) <= 0;
			input_data_tb(636) <= 0;
			input_data_tb(637) <= 0;
			input_data_tb(638) <= 0;
			input_data_tb(639) <= 0;
			input_data_tb(640) <= 0;
			input_data_tb(641) <= 0;
			input_data_tb(642) <= 0;
			input_data_tb(643) <= 0;
			input_data_tb(644) <= 0;
			input_data_tb(645) <= 0;
			input_data_tb(646) <= 0;
			input_data_tb(647) <= 0;
			input_data_tb(648) <= 0;
			input_data_tb(649) <= 0;
			input_data_tb(650) <= 0;
			input_data_tb(651) <= 0;
			input_data_tb(652) <= 0;
			input_data_tb(653) <= 0;
			input_data_tb(654) <= 0;
			input_data_tb(655) <= 0;
			input_data_tb(656) <= 0;
			input_data_tb(657) <= 0;
			input_data_tb(658) <= 0;
			input_data_tb(659) <= 0;
			input_data_tb(660) <= 0;
			input_data_tb(661) <= 0;
			input_data_tb(662) <= 0;
			input_data_tb(663) <= 0;
			input_data_tb(664) <= 0;
			input_data_tb(665) <= 0;
			input_data_tb(666) <= 0;
			input_data_tb(667) <= 0;
			input_data_tb(668) <= 0;
			input_data_tb(669) <= 0;
			input_data_tb(670) <= 0;
			input_data_tb(671) <= 0;
			input_data_tb(672) <= 0;
			input_data_tb(673) <= 0;
			input_data_tb(674) <= 0;
			input_data_tb(675) <= 0;
			input_data_tb(676) <= 0;
			input_data_tb(677) <= 0;
			input_data_tb(678) <= 0;
			input_data_tb(679) <= 0;
			input_data_tb(680) <= 0;
			input_data_tb(681) <= 0;
			input_data_tb(682) <= 0;
			input_data_tb(683) <= 0;
			input_data_tb(684) <= 0;
			input_data_tb(685) <= 0;
			input_data_tb(686) <= 0;
			input_data_tb(687) <= 0;
			input_data_tb(688) <= 0;
			input_data_tb(689) <= 0;
			input_data_tb(690) <= 0;
			input_data_tb(691) <= 0;
			input_data_tb(692) <= 0;
			input_data_tb(693) <= 0;
			input_data_tb(694) <= 0;
			input_data_tb(695) <= 0;
			input_data_tb(696) <= 0;
			input_data_tb(697) <= 0;
			input_data_tb(698) <= 0;
			input_data_tb(699) <= 0;
			input_data_tb(700) <= 0;
			input_data_tb(701) <= 0;
			input_data_tb(702) <= 0;
			input_data_tb(703) <= 0;
			input_data_tb(704) <= 0;
			input_data_tb(705) <= 0;
			input_data_tb(706) <= 0;
			input_data_tb(707) <= 0;
			input_data_tb(708) <= 0;
			input_data_tb(709) <= 0;
			input_data_tb(710) <= 0;
			input_data_tb(711) <= 0;
			input_data_tb(712) <= 0;
			input_data_tb(713) <= 0;
			input_data_tb(714) <= 0;
			input_data_tb(715) <= 0;
			input_data_tb(716) <= 0;
			input_data_tb(717) <= 0;
			input_data_tb(718) <= 0;
			input_data_tb(719) <= 0;
			input_data_tb(720) <= 0;
			input_data_tb(721) <= 0;
			input_data_tb(722) <= 0;
			input_data_tb(723) <= 0;
			input_data_tb(724) <= 0;
			input_data_tb(725) <= 0;
			input_data_tb(726) <= 0;
			input_data_tb(727) <= 0;
			input_data_tb(728) <= 0;
			input_data_tb(729) <= 0;
			input_data_tb(730) <= 0;
			input_data_tb(731) <= 0;
			input_data_tb(732) <= 0;
			input_data_tb(733) <= 0;
			input_data_tb(734) <= 0;
			input_data_tb(735) <= 0;
			input_data_tb(736) <= 0;
			input_data_tb(737) <= 0;
			input_data_tb(738) <= 0;
			input_data_tb(739) <= 0;
			input_data_tb(740) <= 0;
			input_data_tb(741) <= 0;
			input_data_tb(742) <= 0;
			input_data_tb(743) <= 0;
			input_data_tb(744) <= 0;
			input_data_tb(745) <= 0;
			input_data_tb(746) <= 0;
			input_data_tb(747) <= 0;
			input_data_tb(748) <= 0;
			input_data_tb(749) <= 0;
			input_data_tb(750) <= 0;
			input_data_tb(751) <= 0;
			input_data_tb(752) <= 0;
			input_data_tb(753) <= 0;
			input_data_tb(754) <= 0;
			input_data_tb(755) <= 0;
			input_data_tb(756) <= 0;
			input_data_tb(757) <= 0;
			input_data_tb(758) <= 0;
			input_data_tb(759) <= 0;
			input_data_tb(760) <= 0;
			input_data_tb(761) <= 0;
			input_data_tb(762) <= 0;
			input_data_tb(763) <= 0;
			input_data_tb(764) <= 0;
			input_data_tb(765) <= 0;
			input_data_tb(766) <= 0;
			input_data_tb(767) <= 0;
			input_data_tb(768) <= 0;
			input_data_tb(769) <= 0;
			input_data_tb(770) <= 0;
			input_data_tb(771) <= 0;
			input_data_tb(772) <= 0;
			input_data_tb(773) <= 0;
			input_data_tb(774) <= 0;
			input_data_tb(775) <= 0;
			input_data_tb(776) <= 0;
			input_data_tb(777) <= 0;
			input_data_tb(778) <= 0;
			input_data_tb(779) <= 0;
			input_data_tb(780) <= 0;
			input_data_tb(781) <= 0;
			input_data_tb(782) <= 0;
			input_data_tb(783) <= 0;
		wait for 10 ns;
        wait;
    end process;


end behavior;