library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.Types.all;

package vhdl_constants_all_layers_with_bias is


-- Layer 1 Biases
constant LAYER1_BIASES : bias_array_layer1 := (
 -50, -16, -9, -42, -49, -69, -38, -14, -68, -28, -15, -23, -14, 2, -91, -17, -10, -22, -25, -30, -45, -10, -11, -25, -44, 0, -39, 1, -80, 9, 7, 6, -6, -32, -37, -24, 0, -13, -53, 17, -99, -4, 21, -66, -26, 6, -6, -57, -67, 19, -21, -19, -16, 3, -15, -5, 7, -51, -20, 28, -20, -12, -21, 13, 33, -20, -51, 10, -29, -80, 1, -76, -23, -2, -28, -10, 0, 26, -110, -55, -57, -32, -29, 0, 10, -60, -1, -100, -68, -62, -27, 3, -53, -5, -35, -32, -3, 14, -17, 12, -11, 11, 4, -26, -58, -58, -50, -29, 0, -26, -53, 4, 34, -13, -89, -84, -52, -65, -37, 13, -35, -29, -109, 24, -50, 23, -102, 11
);

-- Layer 4 Biases
constant LAYER4_BIASES : bias_array_layer4 := (
 -65, -29, -99, -67, -23, -56, -13, -60, -53, 9, -82, -15, -24, -99, -154, -44, -110, -96, -28, 52, -13, -56, -92, -118, -49, 25, -49, -70, -66, 30, -42, -105, -35, -43, 25, -50, -20, 49, 25, -78, 13, -25, -83, -46, -60, -62, -24, -33, -2, -90, -20, -20, -94, -43, 3, -70, 5, -47, -84, -39, -23, 1, -5, -15
);

-- Layer 6 Biases
constant LAYER6_BIASES : bias_array_layer6 := (
  42, -25, -42, 75, -61, 6, 22, -33, 12, 8
);

end package vhdl_constants_all_layers_with_bias;

package body vhdl_constants_all_layers_with_bias is
end package body;
