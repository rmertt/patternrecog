library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.Types.all;

package Layer4_6_Weights is



constant weight_matrix_layer4 :  weight_matrix_layer4_type := (
  0 => (-37, 79, 40, -65, 7, -43, 87, -15, 11, 1, -37, -23, 6, -12, 81, -82, 15, -132, -31, 77, -45, 42, -74, 11, 26, 32, -3, 9, -17, -10, 29, 72, -18, -29, -51, -122, -3, -26, 24, -10, -10, -61, 74, -78, 93, -31, -42, -57, 96, 54, -80, 32, 55, 7, -28, -59, 6, -77, -2, 48, 71, -29, 53, -38, -14, -9, 5, -35, -6, 1, 16, 42, -17, 56, 9, -61, 33, -19, -131, -3, 26, 21, 19, -8, 83, -17, 9, 10, -94, -61, 2, -86, 28, -13, 65, -121, 0, -15, 28, -73, 2, -7, 34, 18, -51, -76, -2, -32, -13, -55, 10, 9, -151, -17, -15, -32, -73, -81, 61, 11, -28, -13, -68, -70, 11, 2, 29, -6),
  1 => (17, 63, 30, -80, -2, -86, 92, -58, -7, -59, -23, -3, -10, 79, 31, -34, 54, -27, 6, -19, -8, -30, -74, -27, 26, 50, 24, -2, 26, -25, -25, 23, 48, -24, -72, -36, -1, -77, 3, 47, 11, -24, 90, -26, -20, 21, 2, -19, 13, -66, 44, 26, 14, 21, 15, -63, 13, -79, 1, 47, 7, 85, 68, 56, -3, -68, -32, -20, -115, -3, -8, 18, -13, 14, 48, -108, -21, -37, -93, 0, -75, -4, -106, 22, -123, -1, 20, 21, -36, -47, -3, -6, -16, -72, 75, 8, 89, -27, -9, -13, 65, -7, -19, 84, 35, -91, -10, -34, -78, 22, -22, -40, 7, -116, -12, 56, -35, -23, -4, 48, 17, -49, -5, -40, 6, 52, -3, -23),
  2 => (39, 28, -36, -1, 58, 66, 15, 9, -20, 37, 19, 13, 34, 28, -26, -72, 18, 114, 80, 0, -11, 53, 103, 83, 54, -32, 62, 88, 38, -23, -141, -34, 32, 22, 43, 21, -84, -32, -25, 28, -36, -44, 3, -12, -14, -30, -21, -55, -25, -9, -53, -7, 38, -107, -4, 48, 36, 41, 38, 0, -90, 20, 66, -14, 37, 40, 34, -99, -21, 46, 29, 33, -29, 88, 25, 35, -78, -6, -32, -75, -43, -7, 29, 4, -101, 16, 10, -36, 125, 122, -49, -34, -7, 6, -42, -19, 19, 71, 35, 73, 29, 9, 10, 10, 107, 14, -12, 84, -38, 12, -1, 81, -37, -2, 70, -10, 38, 13, 13, 49, 17, 80, 33, 6, -56, 64, 1, -23),
  3 => (10, -47, 0, 73, 16, 50, 35, 85, -10, -41, 11, -15, -7, 63, 17, 55, 29, -34, -58, 19, 36, 2, 15, -72, 12, 12, -38, -7, 82, 52, 38, 12, -47, -4, -34, -47, 55, -70, -72, 11, -9, -32, 31, -14, -1, 85, -84, -8, -42, -80, 33, -49, 46, 16, -95, 16, 60, -6, 4, -21, 37, 3, -42, 66, -78, -41, 56, 39, 16, 7, 6, -21, 74, -35, 6, -17, 41, -88, -17, 14, -42, -5, -4, -66, -22, -59, 49, 27, -3, 1, 6, 35, -50, 19, -5, -46, -27, 32, -31, -29, -24, -93, -8, 8, 28, -46, -24, -16, -109, -35, -35, 80, -28, 55, -31, -41, 90, 26, 6, -29, 1, -86, 52, -60, -94, 5, 98, 30),
  4 => (70, -2, -46, -25, 8, -15, -39, -50, -70, -13, -28, 40, 16, 80, 51, -10, -11, -18, 13, -34, -17, 46, -12, 1, 101, -9, 79, -83, 29, -28, -86, 34, 27, -168, 22, -41, -37, 11, -41, 5, -42, 29, 37, 71, -22, 51, 69, -30, -11, -62, 8, -23, 33, -17, -29, -31, 28, -32, 25, 1, -23, 62, 40, -46, 55, -34, -19, -30, -97, -3, 10, 10, -93, 16, 80, -18, -85, 9, -7, 40, -58, -30, -58, -66, -74, 7, 8, -45, -25, -86, -18, 29, 65, -56, -37, 108, 32, -54, -13, -8, 5, -27, -34, -40, -16, -6, -33, 46, 32, -13, -14, -23, 80, -126, 78, 69, -76, -52, -58, 22, 76, -1, -51, -102, 10, 57, -17, -54),
  5 => (-54, 57, 0, -23, -25, -42, 29, 9, -57, 1, 26, 18, 50, -86, 38, 60, 36, 49, -27, -66, -44, 62, 0, 48, 12, 28, 36, 83, -21, -14, 13, 39, 46, 43, -4, 53, -21, -9, 46, 29, 10, 13, -110, 16, -12, -25, 44, 38, 2, -47, -23, -13, -19, 28, 89, -70, -52, 70, -36, 66, -19, 37, -24, -39, 58, 32, -125, -46, -2, 2, 0, -43, 0, 2, -15, 49, -12, 55, 11, 0, 96, -10, 56, 55, -37, 15, 18, -16, 26, -9, -58, -44, -8, -43, 31, -27, 46, 23, 54, 8, 3, 54, 90, -17, -54, 60, 53, 1, 30, 77, -34, 64, 1, 38, -9, -35, -39, -54, -52, -45, 54, 29, -62, -27, -18, -10, -38, 45),
  6 => (-4, -84, -22, 3, -40, 63, 58, 59, 67, 18, -66, -18, 30, 14, 102, 42, -79, 10, 23, -34, -23, -23, -9, 28, 70, 14, -41, -95, 40, 55, 86, -39, -32, 40, 18, 4, 95, 110, 31, 5, -38, 42, 49, 55, 13, 131, -9, 0, -31, -10, 51, -23, 51, 116, -2, -49, -21, 18, 41, -24, 88, -86, 2, -22, 7, -82, 55, -5, 21, 11, -48, 11, 54, -54, 7, -10, 47, -55, -4, 3, -28, 5, -60, -24, -3, 53, -32, 41, -29, -80, 48, 22, -33, -30, -22, 14, -106, 52, -29, 17, 26, -25, -62, -29, -59, 33, -14, 6, 31, -107, -2, -69, 64, 1, 37, 27, -21, 53, -41, -16, 50, 26, 85, 101, 12, 8, 76, 49),
  7 => (13, -10, 43, 17, 85, 7, -64, -5, -5, 7, 67, 14, 72, 57, -23, 19, 63, -22, -68, -18, 37, 18, 18, -62, 46, -88, -38, -1, 17, 15, 20, 80, -30, 55, 91, -27, -82, 11, -12, 84, 85, 28, 9, -50, 92, -42, -5, 13, -42, 23, -35, -4, 139, 26, 44, 22, -34, -25, -31, -118, 55, -30, -56, -21, 30, 15, 124, -1, -19, -63, -15, -64, -37, -30, 45, 75, -46, 30, 0, 88, -27, -33, -27, -21, 10, -29, -5, -35, 17, -50, -13, 45, -32, 41, -74, 32, -39, 78, 76, -98, -72, 27, 31, 24, -89, -54, -24, 43, -11, -55, -30, -58, -33, 15, -19, 87, 13, -36, -11, 16, 4, -12, 25, -39, -39, -22, 38, -17),
  8 => (35, 11, 47, 14, 9, 54, 7, -61, 10, 4, -97, 29, -17, -27, 46, -64, -112, -14, 39, 25, -87, 45, 25, 28, 68, -68, 13, 52, -25, 18, 3, 28, -7, -34, 47, -38, -32, 21, 73, -76, 7, -12, -45, 59, -25, 30, 15, 22, 10, -57, -52, -2, -32, 34, 1, -29, -26, -53, -22, -16, 34, -33, 2, -112, 39, 21, -2, 23, -65, 2, -68, 5, -169, 13, -52, -35, 33, 37, 33, 33, -17, -7, -127, -28, -32, 60, -89, 9, 13, -16, 16, -115, 35, 59, -22, 23, -37, -20, 76, 23, -27, 13, -23, 19, -8, -69, 82, 45, 36, -18, 4, -112, -20, -109, 59, 96, -79, -71, -18, -5, 12, 22, -16, -59, 1, -49, 18, 31),
  9 => (0, 2, 30, 111, 17, 42, -8, -31, 59, -62, -47, 48, 28, 102, 34, -66, -20, -37, -26, -77, -44, 34, -29, 3, 83, -95, 75, 45, 2, 42, 48, 3, -23, -83, 13, -40, 103, -62, -69, -44, -50, -48, 95, 44, 0, 2, -50, -76, 67, -22, -72, -30, -16, 40, -12, 32, 36, -70, -8, 7, 102, 33, 41, 27, 8, 11, 58, 44, -89, 81, 45, 131, -150, -72, 45, -32, 54, -36, 21, -58, -3, 5, -43, 9, 13, -81, -59, -41, 73, -57, -28, -47, 22, 89, 23, 7, -37, 29, 69, -7, -42, -21, -97, 22, 62, -53, -12, 34, -55, 16, 46, -20, -25, -56, 76, 10, 21, 12, 5, 69, 35, -6, -14, 2, 13, 53, 86, -65),
  10 => (3, -29, 3, -8, 10, 41, 36, 58, 54, 23, 3, -1, 71, 0, 11, 42, -3, 69, -2, -18, 2, 24, -7, 35, 31, 29, -65, 8, 34, 30, 42, -32, -31, 77, -11, -9, -5, 30, 64, 40, -55, 20, 36, 33, -41, 55, 30, 56, 28, 7, 70, -16, 58, 72, 19, -87, 23, 34, 61, -37, 17, 20, 16, -2, 2, -35, 39, -15, 84, -40, 26, -50, 44, -117, 11, 49, -36, -2, -14, 48, -3, 28, 21, -23, 1, 26, -9, -15, -51, -141, 12, 45, 28, -86, -2, 51, -26, 86, -76, 52, 4, 24, -2, 1, -60, 95, -6, -11, -21, -53, -20, -8, 122, 40, 10, -9, 10, 84, -35, -2, 133, 48, 79, 154, -46, 45, 31, 40),
  11 => (-57, 36, 14, -5, -83, 38, -56, -45, -39, 67, -64, -18, 9, 34, -94, 67, 0, -4, -150, -51, 26, 5, -19, 15, 13, 57, 47, -31, 0, 55, -4, 9, -38, 62, -79, -48, -20, -37, 54, -12, 42, 41, -39, 39, -29, -5, 16, -12, 31, 76, 7, 21, -81, 40, 46, -10, -82, 52, -11, 47, -32, 98, -25, 68, 28, -51, -106, 21, -11, 56, 96, -56, 40, 15, -15, -9, -2, -95, 51, -56, -26, -77, 65, 10, -33, 6, 41, 10, -14, -75, -11, 100, -39, -68, 32, -53, 53, -61, 17, -41, -13, -31, 38, 45, 17, -68, -59, -89, -4, 158, -80, -41, -18, -69, -60, -45, -27, 102, -74, 46, -13, -35, -4, -6, -23, -32, 0, -8),
  12 => (17, 52, 94, -13, -47, -124, -60, -45, 101, -18, -32, -5, 151, -13, -27, 41, 54, 35, 15, -39, -30, 119, 84, 50, 45, -90, -65, 97, -36, 18, 63, -9, -13, 22, -17, -1, 12, -20, 1, -64, 74, -2, 18, 41, 9, -106, -33, 74, 81, -75, -52, -90, -43, 19, 31, -10, -94, 0, -65, 25, -12, 73, 31, -46, -68, -24, -19, 24, -50, -22, 48, -46, 27, 10, -40, -105, 48, 9, -3, 9, 9, -50, 40, -21, -25, -7, -104, 15, -10, -44, 103, -9, 7, -1, 52, -55, 43, 34, -15, 13, -78, 4, 23, 19, 11, 18, 50, 46, 71, 8, 49, 38, -46, -39, -13, 3, -72, -41, 71, 6, 22, 89, -25, 54, 27, -22, -31, -68),
  13 => (105, 23, -7, -6, -14, -14, -106, 49, -8, -3, 8, -18, -53, -7, -55, 10, -62, -13, 62, 6, 32, -50, 32, 18, -4, 54, -23, -24, -20, 52, -2, 11, 56, 14, 97, -7, 2, -24, -28, 25, -7, 61, -10, 3, 5, -2, 57, 31, -4, 34, 54, -11, 4, -9, -118, 78, 43, 49, 62, -6, -3, -8, 94, 55, -31, 8, -2, -17, 49, -6, 13, -84, 22, 10, 32, 34, -49, 45, -53, 6, 50, 19, 19, -67, -49, -51, 51, -48, 83, -9, 32, -42, -48, -73, -56, 46, -56, 59, -51, 58, 32, 93, -31, 36, 29, 21, 72, 105, 43, -13, 98, 95, 73, 11, 64, -19, -9, 11, 93, -4, 43, 28, -4, 39, 69, 54, 23, -30),
  14 => (44, -42, -36, -41, -45, -32, -72, 19, 2, 122, -77, -41, -11, 4, 19, 59, -55, 64, 70, 86, -68, -23, 23, 3, -19, -2, 20, -71, -27, 57, -17, 35, 51, 52, -32, -58, 14, 21, 24, -27, 8, -9, 31, 55, 71, -29, -12, 58, 48, 39, 59, 59, -27, 50, -13, 66, -41, 109, 9, 29, -1, -75, 83, 33, 89, 17, 28, 55, 39, 109, 19, 4, -2, -4, -7, -12, 3, 19, 12, 28, 47, 21, -28, -5, 14, 75, -3, -30, -45, -63, 44, 23, -36, -26, 66, -70, 60, -1, 42, -58, 14, 46, 8, -34, -3, 23, 85, 122, 59, 77, 40, -24, 14, -44, 18, -51, -2, 49, -12, -13, 59, 74, 62, -16, 72, 2, -22, -27),
  15 => (-36, 143, 26, 69, -21, 41, -47, -85, -33, 40, 51, 12, -13, -86, -11, 52, 34, -49, -107, -52, -10, -15, 13, -86, 10, 34, 50, -59, 21, 16, 22, -76, -69, 44, -43, 8, 23, 8, 19, -6, -68, 10, -31, -34, -88, 18, -7, -12, 47, 19, 78, -3, -33, -37, -35, -37, -16, -72, 15, -67, -57, 151, -41, -6, -14, -54, 1, 54, 9, 33, 63, -32, 16, -26, 22, 32, -23, -16, 72, -28, -40, -30, -82, -64, 15, 4, -7, 30, -33, -25, -2, 53, -64, 24, 32, -31, 88, -3, -58, -123, -79, -39, 3, 38, -31, -34, -56, -124, -74, 101, -108, -57, 15, -21, -88, -17, -47, 48, -57, 104, -38, -100, 19, -22, -71, -25, -14, 52),
  16 => (-19, 75, 92, -27, -47, 26, 66, -50, 25, -52, -49, -36, 51, 35, 5, -5, 14, 28, -24, 11, 13, 60, 33, -33, 95, -34, 35, 6, 8, -44, -31, 47, -80, -74, -73, -52, 9, -46, 4, 44, -14, -25, -5, 5, -28, 87, -7, 18, 32, -43, 44, -79, -22, 77, 16, -91, 40, -55, 68, -68, -27, 81, 31, -15, -23, -44, -23, 27, -110, -40, -9, 27, -66, -34, 75, -43, -96, -98, -3, -1, -73, -48, -23, -25, -64, -49, -20, 30, -21, -19, 0, 53, 48, -72, -15, -14, 53, 29, -36, -7, -38, -34, -33, 105, -29, 18, 6, -59, -21, 36, -68, 29, 51, -60, -20, 32, -26, -9, -9, 91, 10, 6, -1, -110, -24, 53, -35, 4),
  17 => (18, -47, 81, -30, -11, -109, -44, 81, 110, 11, 43, 6, 95, 41, -51, -30, 0, -39, 22, 47, 74, 67, 18, 20, 40, -80, -76, 36, 95, -41, 43, -52, -27, 93, 62, -8, -34, -103, -77, 30, 35, -35, 67, 22, -12, -129, -8, 13, 4, -22, -88, -46, 32, -6, 43, 58, 16, -24, -100, -135, 34, 30, 8, -8, -8, 1, 62, 28, 51, -128, -1, -80, 17, -63, 39, -31, 24, 2, -11, 46, -51, -44, -42, -75, -54, -33, -13, 1, -25, -45, 91, 4, 15, -17, -42, 4, -46, 43, -8, -44, -15, 17, 38, 58, -1, 33, -44, -3, -32, 37, 11, -31, -65, -15, 50, 40, 73, -74, 27, 32, -26, 56, -19, 12, -71, 1, -41, -30),
  18 => (-2, 103, -13, 21, -2, -31, 12, -31, -124, 49, -38, -19, -1, -90, 37, -9, -15, 50, -103, -20, -72, 37, -59, -16, -33, 57, 63, 49, 6, 13, 3, 84, -15, -15, -60, -3, 34, -32, 58, 70, -34, 14, 16, -48, 59, -47, -17, 33, 23, 7, 49, -59, 48, -35, -37, -61, 2, 54, -23, 71, 10, 107, 57, 46, 34, -13, -61, 84, -9, 56, -57, 93, -33, -3, 49, 9, 45, 8, 107, -13, 47, 38, 85, 49, -20, -73, 39, 5, 19, 50, -65, 18, -4, 92, -5, 33, 66, -68, 59, -20, -22, -31, 26, -57, 37, 6, 34, -69, -4, 86, -41, 63, 10, 81, -53, -21, 11, 36, 10, 75, 8, -57, -143, -71, 9, -4, 14, -35),
  19 => (72, 26, 47, -20, -92, -15, -86, -4, -8, -93, -47, -50, 82, -79, -26, 99, -7, -20, -21, -69, 41, 77, 55, -1, 65, -65, -63, 45, -38, 23, -10, 3, -58, 47, -15, 13, 15, -98, 31, -85, 35, 54, -86, 3, 2, 9, 0, 107, 42, -65, 61, -98, -64, -1, 45, 27, -93, 47, -17, -47, -23, -12, 48, -73, -79, 21, -85, -27, -63, -29, 58, -35, 1, 53, -41, -4, -1, -59, 32, 83, -8, -96, -1, -49, 29, 7, -112, 2, 23, -45, 62, -9, -25, -33, -43, 53, 23, 18, -26, -100, -126, -13, 24, 28, -33, 48, 16, -18, 50, 32, -15, 79, -53, -50, -21, 27, -32, -12, -49, -80, 72, 2, -38, 17, 39, -81, 11, -23),
  20 => (75, -4, -40, -8, 44, -82, 13, 49, 36, 16, 65, 54, 3, 47, 41, 85, 61, -37, 21, -28, 51, -44, -44, -98, -30, -38, 17, -61, 40, -75, -24, 99, 43, 62, 84, 12, -20, 62, 33, -9, 9, 83, -2, 7, 38, -102, 28, -17, -37, 52, 54, 86, 60, 19, 2, 24, 36, 57, -49, 2, -42, 17, -129, 22, 41, 37, -27, 99, 107, 38, 79, 82, -25, -38, -10, 100, -21, 86, 59, 50, 7, -30, -69, 66, 56, -19, -6, -54, -55, 22, -29, 39, 35, 7, -65, 22, 38, -52, 47, -31, 39, 46, 17, 12, -87, 40, 13, 15, 51, 16, -84, -1, -13, 25, 17, 90, -8, 65, 7, -19, 49, -37, -21, 82, -4, -7, -62, -83),
  21 => (-89, -7, -14, -47, 23, -21, 16, -9, 23, -13, 77, 42, 29, -83, 41, 81, 15, -83, -14, -9, 59, -11, -45, -44, -20, 43, -83, -62, 30, -3, 80, 6, 49, 52, 51, -47, 68, -16, 58, 18, -23, -15, -44, -74, -20, 15, -27, 53, -2, 39, 85, 40, -30, 77, -23, 4, 40, 30, -37, 2, 39, 42, -53, 21, -77, -29, 40, 73, 65, 3, 44, -40, 79, 8, -55, 79, -16, 41, 8, -82, 82, -39, -18, 34, 34, -46, 29, -39, -62, 2, -49, 28, 11, -43, 27, -64, -18, -25, -3, -81, -10, 47, 16, -5, -123, 105, -6, -5, 42, -12, 0, 35, 74, 11, -37, -16, 3, 29, -23, -39, 26, -3, 25, 18, 18, -41, 10, 23),
  22 => (-86, 27, 48, 23, -8, 12, -50, 30, 80, -34, -12, 14, 65, -21, 5, 7, 29, -20, 22, 81, 62, 51, -21, 31, 80, -28, 18, 44, 1, -53, 5, -2, 17, 4, -23, -84, -39, -58, -54, 14, 3, -153, 56, -57, 2, 21, -138, -46, 6, -9, -25, -23, 78, -8, 49, 33, 99, -24, 35, -49, -19, 28, 39, 24, -75, 33, 34, -39, -42, 22, 30, 16, -2, 68, -15, -72, 16, -25, -21, -70, -54, -37, 18, -139, 1, 2, 52, -54, -1, 29, 63, 14, -33, -17, 46, -129, 49, 43, 5, -88, -33, -24, 16, 56, 3, -23, -33, -10, -64, 16, 23, -9, -78, -33, -34, -81, 9, -6, 40, 55, -66, 15, 8, -53, -53, 36, 14, -1),
  23 => (-5, 44, 7, 26, 3, 53, 18, 13, -42, 5, -1, 3, -23, -18, 24, 12, -26, 83, -30, 41, 30, -31, -56, 24, -9, 67, -10, -7, -21, 66, -14, -11, -58, 11, -73, 2, 20, 91, 17, -44, -4, 4, 54, 65, -70, 22, 3, -48, 99, -31, 31, 44, -57, -23, 49, -59, 71, 59, 42, 1, 34, 6, 4, -55, -54, -28, -20, -94, 33, -58, -86, -52, 57, -70, 90, 6, 17, -24, -107, -45, 25, 50, 22, 48, -11, 3, -5, 37, 37, -16, -23, 21, -4, -15, 54, -12, -5, -4, -60, 46, 36, -48, -12, -12, 8, 7, -19, -7, 9, -3, 8, 41, 50, 46, -12, -23, -22, 34, -8, 16, 18, 22, 83, 62, -6, -15, 95, 85),
  24 => (33, 2, 35, -56, 25, 46, 5, 68, -64, 1, 34, 48, 54, 34, -2, -23, 91, 12, -37, 3, -19, 45, 16, 3, 6, 32, -79, 35, 50, 47, -69, 11, -68, 83, 2, 81, -41, 17, 23, 52, -5, -9, -51, -30, 26, 23, -27, -55, -16, -14, -38, -25, 31, 10, 80, 2, -12, 56, 72, -30, 66, -17, -122, 33, 29, 40, 28, -33, 61, -58, 41, 44, -16, -71, 49, 62, -27, 6, 11, -13, -34, 13, -36, 38, 3, 26, -24, -78, -93, 52, 6, 39, 47, 1, -30, 19, 85, 87, 32, -23, -97, 14, 53, 34, -11, 55, 19, -56, -23, 46, -18, 34, 15, 18, -61, 28, -2, -28, -12, 48, -45, -83, 60, -67, -72, 4, 57, 60),
  25 => (7, -2, -10, -41, -23, 11, -23, -4, 1, 50, -51, 23, -14, -3, 23, 128, 30, 3, -30, 41, -5, -4, 31, -119, 10, -25, 6, 10, 7, 61, 93, 68, -46, 40, -3, 24, 95, -11, 14, -2, -7, -7, 19, -66, 56, 0, -48, -52, -28, 12, 98, 30, 52, 49, -8, 64, 42, 76, 44, -8, -36, 2, -10, 69, -46, 52, 27, 74, 87, 17, 29, 32, 57, 13, -80, 0, 17, -89, 36, 19, -8, -18, 8, -16, 52, 52, 24, 26, -5, -6, -8, 76, -39, 16, 35, -44, 23, -40, -51, -130, -19, -44, 38, -41, -3, 29, -5, -5, 15, 51, -35, -22, 43, 104, -81, -35, 111, 151, -65, -7, -30, -7, 64, 41, -44, -23, 36, 8),
  26 => (54, -46, -11, 53, 37, 66, -46, 34, -52, -51, 47, -41, -14, -25, -43, 22, -95, -60, 34, -38, 67, 11, -1, -7, -54, 32, 0, -30, 60, 102, -15, -7, -8, -64, 26, -43, -40, -37, -10, 75, -41, 88, 105, 1, -30, 0, 67, 15, 3, -37, -39, -15, 20, 3, -29, -110, 60, 20, 62, -40, -8, 60, 18, 3, 12, -46, -20, -45, -46, -62, -17, -57, 32, -24, 63, 69, 14, 56, 9, -27, -1, 65, 15, -57, -20, -60, 5, -10, -31, -57, -81, 10, 56, 7, -20, 103, -25, 9, -94, -12, 7, 21, -51, -68, -39, 15, 32, -20, 2, -22, 25, 59, 34, -61, 110, 48, -101, -55, 34, 15, 90, -32, -19, 10, 4, 81, -15, 46),
  27 => (9, 23, -55, 146, 46, 90, 36, -69, 24, -15, -24, -29, -13, 24, 29, -13, -45, 78, 31, -11, 10, 23, 58, -14, 72, -32, 109, -46, -29, -20, -7, 59, -4, 7, -28, -9, 33, -92, -2, -82, 61, -44, 9, 22, 40, 74, -8, 3, 15, -69, -2, -7, 0, 16, -77, 20, -33, 57, -20, -13, 3, 7, 108, 24, -24, -7, 31, 20, -60, 80, -18, -10, -37, 28, -45, -69, 22, 10, 28, 27, -69, -55, -9, -56, -55, 21, -37, 53, 96, 74, -4, -11, 40, 93, -43, -41, 58, -22, 21, 82, 47, -25, -85, 46, 57, -73, -19, 0, -27, 12, 16, 37, -40, -65, 36, -25, 35, -29, 26, 46, -6, 4, 18, -63, 42, 29, 97, 41),
  28 => (45, 19, -16, -99, -49, -101, -62, -51, 100, 76, 56, 43, 49, 83, -10, 59, 36, 46, 24, 62, -37, -11, 48, 16, -26, -46, 43, 19, 6, 1, -49, 4, 13, 42, -2, 54, -49, 128, -15, -7, -7, 35, -4, 47, 23, -120, 21, 48, 3, 59, 45, 30, -45, 4, 31, 81, 41, 35, 22, 20, -50, -7, -77, 37, 25, 49, 35, 20, 83, 107, 38, 31, -20, -39, 48, -6, -42, 19, 36, 8, -37, -26, -23, -64, 33, 23, -1, -86, -35, 39, 79, 62, 0, -26, -29, 39, 42, -19, 11, 35, 60, 27, 10, 17, -27, -16, 31, 88, 41, 63, 32, -25, 27, 31, 30, 17, 80, 117, -21, 29, -8, 82, -16, 126, -35, 61, -101, -99),
  29 => (-56, 36, -44, -70, 28, -22, 44, -1, 56, -28, 76, 85, -57, 33, 67, -43, 18, -92, 2, -9, 127, -6, -72, -3, -51, 51, -62, -34, 46, -138, -11, 15, 10, -43, 39, -38, 37, -12, 11, 126, -69, -30, 15, -12, 24, -12, -8, 0, -23, 40, -23, -31, 64, 93, -41, 5, 120, 11, 38, -74, 52, 28, 22, 43, -101, -46, 10, 27, -16, -48, -63, 57, -3, -113, 72, 68, 36, 75, -40, -28, 29, -28, -20, -8, 39, -61, 63, -42, -117, 9, -43, -14, 48, -37, -49, -4, -26, 2, -1, -106, 18, 46, -30, 25, -69, 40, 25, 39, 20, -29, 47, -85, -4, 18, -21, 0, 19, -14, 57, -39, -32, -26, -8, 8, -14, 31, 31, 26),
  30 => (57, 96, -15, 27, -96, -10, 39, -52, -44, 15, -125, -91, -65, 30, 43, 12, 23, 13, -63, -55, -97, 8, -69, 15, 36, 55, 90, -8, -18, 44, 17, 11, -65, -75, -115, 26, -31, -44, 5, -89, 58, 19, 31, 57, 31, -25, -3, -33, 75, 1, 63, 50, -80, 24, 31, -35, -4, 9, -43, 94, 25, 34, 21, -40, -17, 54, -45, -23, -50, 32, 7, 32, -21, -6, 9, -42, 12, -124, 11, 28, -31, -48, 55, 34, 37, 24, -8, 47, -43, 14, -55, 1, -21, -16, 37, -5, 64, -78, 21, 13, -6, -76, 33, 39, 7, -76, 4, -61, -57, 48, -8, 33, -8, 1, -45, -16, 0, -2, -27, 1, 34, -65, -36, -62, -12, -51, 26, -37),
  31 => (-28, -66, 25, 41, -11, 88, -103, 18, 8, -57, 14, 29, 1, 23, -11, -82, 60, -104, -96, 25, -18, 85, -15, -49, 28, -77, -1, -45, 16, -32, 28, -37, -6, 36, -45, -41, 10, 29, -2, 10, -4, -21, 58, -21, 26, -4, -6, -15, 115, 18, -122, -33, 17, -56, -65, -43, 47, 32, 5, -20, -44, 97, -56, 10, -31, -7, -18, -59, 21, -13, 23, -61, 54, -85, 60, -10, 26, -35, 102, -12, -10, -2, 4, -39, 103, -56, -13, -84, -46, 17, -19, 22, 15, -3, 85, 23, -47, 14, 20, -19, 25, -58, -4, 100, -104, -1, -39, -124, -31, 48, 2, -8, -15, 46, -10, -12, 16, -73, -35, -3, -15, 3, 9, -8, -52, -24, 2, 94),
  32 => (88, 33, -63, 5, -41, 15, 9, -82, -91, 31, -88, -37, -57, -49, 36, 40, -64, -86, -67, -47, -61, 0, -60, -28, -54, 27, -8, -6, -18, 75, 15, 17, -25, 51, -34, 69, -4, -38, 69, -34, 38, 103, 19, -20, 37, 5, 34, 47, 59, -15, 62, 55, -66, -1, -31, -87, -90, 50, -57, 6, 9, 30, 36, -63, 34, 16, -17, 17, 15, 8, 8, 40, -1, 2, -15, 5, 42, -10, 71, 85, 5, 6, 64, 48, 40, 86, -34, -26, -38, 18, -29, -12, -19, 56, -6, 21, 13, -97, -8, 7, -88, -40, 33, 1, 32, -45, 30, -29, -41, 28, -6, 59, 52, 16, -49, 30, -48, 20, -1, 37, -6, -33, -94, -59, 33, -80, -39, -28),
  33 => (-78, 27, 11, 48, 54, 44, -23, -40, 8, 26, 8, 29, -8, -44, -2, -18, -19, 17, -52, -38, -25, 17, 20, 16, 1, -16, 63, 48, 47, -75, 1, 23, 31, -79, -17, -25, 32, -70, 11, -66, 59, -107, -50, -99, 61, 44, -71, -8, 40, 0, -23, 8, 29, -11, 4, 11, -18, 18, -38, -63, 34, -8, -12, -8, -17, 55, 19, 16, -77, 55, 35, -21, -36, 66, -37, -81, 102, -33, 85, -38, -5, -115, 68, -19, 62, 22, 62, 60, 100, 42, -25, -19, -22, 67, 12, -86, -10, -19, 67, -26, 20, 9, -7, 4, -15, -28, 20, 26, -18, 60, -12, -80, -107, -54, -85, -92, -21, -26, -59, 32, -76, 12, 21, -107, 13, 19, 29, 62),
  34 => (93, -14, 39, -58, -35, -44, -30, 9, -45, -53, 28, -41, 37, -48, -6, -43, 8, 3, -44, -15, 40, 33, 9, 8, 18, -31, 10, -15, -2, 9, 25, 79, 15, 16, 54, 11, 9, -53, 92, 5, 9, 80, -30, 78, 26, -5, 118, 23, 17, 27, -70, -62, -29, -8, 19, -5, -34, -7, -111, -30, -31, 26, 50, -48, 29, 39, -43, 24, 21, -44, -46, 8, 29, -7, 32, 44, 2, -12, 88, 36, 49, -19, 7, -6, 46, 49, -4, -4, 2, 27, -32, -71, 99, -64, -32, 104, 7, -55, 18, 26, -60, -30, 15, 41, -85, -17, 26, 14, 40, 2, -31, -9, -46, 19, 43, 113, -67, -96, -16, -31, 88, 13, -103, 46, 83, -48, -40, 14),
  35 => (-1, -86, 22, 18, 77, 27, -51, 7, 7, 34, 9, 64, 29, 41, -31, -47, -92, 54, 113, 19, -4, -1, 66, 14, 41, -18, 48, 5, -6, 23, -50, -12, 154, 75, 106, -41, -19, 27, 5, 15, -11, 11, -9, 32, -31, -46, 5, 10, -29, 33, -82, 9, 35, -29, -13, 58, 38, -44, 21, -14, -61, -58, 16, -3, 29, -15, 61, -63, -39, 64, 8, -31, -24, 61, 13, -28, -47, 147, -45, -2, 36, -25, -32, -50, -40, 13, 80, -33, 37, 43, -6, -100, -1, -27, -75, -19, -48, 0, -11, 43, 42, 140, 20, -13, 15, 17, 69, 105, 110, -39, 75, 32, 2, -100, 105, 64, -48, -23, 64, -24, 1, 45, -32, 27, 78, 23, -9, -37),
  36 => (113, 23, 14, -59, -105, -55, -64, 17, -23, -13, -76, -55, 46, -10, -31, 15, -13, 12, -27, -30, -82, 18, -47, 77, 3, 8, 50, 12, -70, 53, -21, -28, 22, 33, -5, 72, -2, 54, 32, -55, -8, 80, 16, 106, -33, -92, 115, 67, 37, 7, 42, -2, -63, -36, 60, -56, -67, 42, -30, 48, -64, 26, 42, -28, 42, 5, -89, -37, 11, 1, 26, -75, -8, -22, 31, 4, -55, -3, -7, 84, 69, -39, 43, 83, -13, 79, 27, -25, -27, -31, 10, 41, -13, -71, 25, 64, 37, 18, -58, 92, 25, 34, 21, 5, -34, 17, 51, -5, 55, 55, 12, 34, 34, -41, 55, 70, -100, 10, -31, -16, 70, 25, -59, 46, 44, -86, -50, -81),
  37 => (36, -75, -54, 0, 25, 17, 37, -12, -12, -58, 11, 63, -42, 8, 42, -71, -46, -9, 16, -58, -15, -16, -48, 47, -16, 45, 2, -79, 68, -88, 10, -1, 30, -16, 36, 23, 50, 10, 65, 15, 62, 24, -49, 10, 34, 64, 23, 43, -65, 14, -86, -57, 4, 35, -43, -45, -44, -44, -127, 42, -14, -13, -58, -69, -59, -19, 27, 35, -7, 1, 9, -8, -18, 12, 35, -57, 46, 42, 8, -6, 39, -65, -44, 29, 37, 59, 8, 9, -7, 42, -24, -22, 75, 18, -49, 58, -48, -82, -26, -23, 25, 45, 55, -41, -65, -22, 27, 30, 47, -87, -38, -52, -33, 3, -47, 25, -30, -82, -44, -37, -50, -28, -8, -26, -6, -30, 17, -2),
  38 => (37, -49, 6, 21, -23, -3, 47, -53, 58, -7, -70, -4, 59, -62, 20, -14, -36, 16, 19, -41, -61, 81, 62, 54, 63, -56, 126, 33, -53, -84, -17, 35, -17, -36, 25, 30, -52, 25, 46, -109, 82, 36, -38, 86, -41, 8, -34, 67, 19, -16, 10, -30, -59, -7, 61, -37, -59, 38, -34, 11, -37, -40, 5, -141, 37, 9, 4, 0, -18, 104, 1, -34, 16, -3, -127, -40, 26, 7, 53, 76, 35, -75, 16, 47, 0, 44, -99, 28, 19, -42, 26, -75, 53, 3, 9, 33, -10, -20, 64, 42, -3, 25, 26, -4, 0, 42, 47, 18, -13, -30, 5, -106, 3, -50, 16, 5, -56, -14, -141, -21, 57, 2, 38, 12, -12, -73, -25, 60),
  39 => (18, -48, -65, -5, 1, 3, 46, 52, -3, -41, 11, 28, -73, 28, 43, 52, -41, -96, -9, -11, 24, -52, 14, -107, -16, 1, -4, -68, 61, 10, 44, 112, -22, 29, 66, -1, 67, -37, 22, 40, -5, 36, -12, 27, 56, 0, 53, -18, -19, -18, 73, 22, -35, 96, -46, -19, 44, 24, -30, -52, 43, -1, -96, 26, -22, 32, 47, 146, 54, 20, -45, 69, 6, -84, 8, 70, 66, 27, 52, 19, 9, -21, -84, -6, 39, 6, 23, -11, -43, -15, -30, 26, 50, 32, -85, 54, -23, -49, 40, 13, -6, 58, -52, -10, -55, 18, 4, 35, -30, -60, -8, -32, 37, 52, -22, 40, 68, 63, -51, -28, -5, -6, 77, 26, -58, 43, -6, 25),
  40 => (-16, -4, 55, 47, 82, 52, 11, 63, -50, -78, 72, 9, 34, 49, 95, 5, 16, -89, -61, -61, 104, 32, 20, -83, 54, -17, -64, 41, 108, 2, 30, 56, -84, -36, -21, -32, 59, -59, -79, 120, -74, 5, 8, 10, -65, 35, -47, -57, -29, -19, 33, 5, 83, -44, -90, -48, 18, -53, 13, -13, -1, 23, -15, 61, 1, -50, -2, 14, -91, 27, 16, -1, 66, -14, -6, 59, 23, -41, -5, -63, -33, 9, -18, -44, -22, -21, 43, -24, -46, 21, 16, 22, 16, 45, -36, -18, 37, 24, -7, -82, -8, -9, 41, 16, 12, -31, -66, 14, -99, -40, -68, 6, -47, -25, -124, 2, 23, 51, -63, -15, -31, -59, -20, -22, -83, 54, 27, 20),
  41 => (-142, 26, -1, 34, 128, 31, 10, -41, 3, -39, 85, 131, 5, 61, -21, -24, 17, 24, 24, 13, 16, -9, 19, -22, 5, 50, 43, 46, 1, -60, 13, -47, 78, 12, 62, -69, -12, 79, -82, 52, 6, -111, 96, -109, -39, 23, -111, -55, 44, -12, -44, 3, 45, -70, -18, 73, 70, 4, 68, 6, -7, 54, 14, -3, -68, 19, 48, -35, -58, 44, 67, -19, 28, 19, 11, -5, 27, 17, -33, -127, -19, -18, -47, -28, -11, -36, 62, 75, -30, -5, 40, 69, -89, 11, 77, -76, -7, 35, -34, -28, 37, 29, 0, -13, 66, -19, -58, -26, -52, 55, -58, -57, -2, -41, -44, -44, -28, 11, -28, 17, -96, -9, 33, -133, -38, 97, 39, -29),
  42 => (0, -67, -36, 70, -45, 30, 20, 26, 17, 48, -75, 18, -7, 2, -28, 23, -103, 8, 130, 94, -38, -70, 39, 38, -62, -23, 18, -39, -90, -24, 41, 54, 62, 34, -35, 43, 38, 32, -32, -79, -29, 9, -9, -13, 51, 41, -16, 30, -28, 19, 24, 25, -31, 74, -54, 45, 13, 40, 20, -48, 89, -70, 38, 8, 12, -25, 24, 66, 45, -15, -50, -46, 10, 66, -76, -34, -5, 84, -13, 20, 63, -21, -47, -41, 40, 37, 21, 7, 15, -26, 40, -63, -92, -63, -30, -46, -24, -2, -17, 32, 17, 73, -85, -31, -34, 46, 89, 99, -6, -32, 95, 28, -13, 15, 105, -50, -12, -31, 108, -23, 40, 62, 2, 18, 71, 0, 40, 76),
  43 => (36, 94, -52, 30, -17, -6, 36, -48, -60, 80, -4, -29, -4, -83, -10, 42, 53, 46, 6, 36, 5, -43, -49, 35, -80, 67, 78, 13, -92, 38, -24, -7, 10, 76, -9, 37, -48, -28, -14, -9, -17, 46, -18, -27, -50, 8, 16, 33, -9, 55, 13, 88, 4, -34, 34, 50, 30, 75, 19, 93, 10, 90, 74, 25, 48, -41, -44, 46, 48, 13, -31, 6, 51, -14, 25, 5, -60, -24, -23, -22, 10, 54, 75, 59, -123, -18, 78, 12, 54, 14, -102, 46, -28, 28, -10, 6, 89, 34, 21, 15, 43, 12, -70, -72, 69, -14, -9, 29, -52, 84, -50, 41, 25, 42, 30, -11, -9, 3, 54, 62, 47, -6, 1, 15, -39, 25, -56, 8),
  44 => (-39, 26, -75, -7, 21, 15, -18, -121, -19, 11, 16, 56, -101, -48, -29, 26, -11, -20, -12, 45, -23, -54, -15, -15, -6, 57, 65, -27, 5, -64, -20, 34, 89, -10, -1, -14, -66, 46, -13, -12, -13, 13, 12, -53, 4, -15, -36, -27, 37, 90, -25, 92, 24, -19, -19, -60, 18, -5, -107, 99, 17, 32, -8, -3, 10, -78, -22, 2, -64, 35, 14, -10, -13, 19, 24, -9, -21, 22, 2, -90, -17, -29, -46, 65, -12, -12, 106, 8, -6, -16, -111, -23, 41, -5, 48, -46, 1, -130, -28, -42, 43, 29, 10, -27, -48, -52, 30, -3, 38, 21, 11, -90, 8, -90, 30, 0, -85, -72, -6, 23, -16, -50, -75, -76, 58, -49, -22, 18),
  45 => (-44, 5, 28, -43, 9, 35, 19, -92, 73, -33, 7, 45, 32, 18, 2, -99, 3, -5, 96, 75, -28, 59, 84, 58, 80, -100, 54, 13, 58, -92, -89, 5, 27, -50, -1, -36, 15, 36, 7, 20, -42, -62, -25, -8, -39, 54, -50, 3, 14, -100, -42, -46, 2, -57, 1, 47, -11, -52, 64, -119, -52, -21, 38, -84, -6, 10, 76, -63, -35, 25, -1, 51, -64, 49, 19, -37, -48, 53, -19, -65, 6, -53, -88, -3, 25, 42, 10, 23, -48, 41, 51, -46, 6, -22, 16, -43, 17, 57, 51, 18, 25, -35, -4, 49, -25, -6, 11, 3, -13, 11, 32, -49, -58, -37, -16, 74, 40, 6, -1, 1, -51, 96, 21, -15, -13, 2, -61, 13),
  46 => (84, -39, 9, 17, 13, 8, 31, -39, -9, -41, -98, 90, 1, 38, 73, -67, -71, -5, -24, 43, -23, 24, -9, 14, 24, -15, -8, 15, 42, 3, 30, -16, -30, -27, 85, -47, 9, 28, 30, -30, 7, 48, -35, 76, 23, 35, 36, -30, -6, -62, -46, -27, -28, 23, 14, -42, -50, -56, -96, -26, 11, -62, 9, -83, 11, -34, 30, -37, 73, 46, -82, 57, -38, -4, -28, 41, 54, 14, 32, 34, -21, -9, -137, -26, 27, 54, -34, 23, 47, -24, -10, -73, 85, 32, -25, 11, -47, -53, 84, 33, -18, -2, 15, -10, -20, -72, 21, 2, 35, -61, 31, -117, -100, -1, 33, 59, 5, -57, -28, -8, 17, -13, 66, -42, -29, -81, 2, 30),
  47 => (-57, -38, -7, 62, 53, 12, 27, 1, -6, 57, -59, 12, -28, 20, 21, 5, 35, -35, 27, -45, -68, -71, -47, 6, 8, -41, 4, -21, 73, -35, 50, 35, 73, 57, 51, 5, 73, -18, 4, -28, 4, -53, -17, -62, 44, 31, -71, -26, -52, 5, -50, 39, 26, 8, 24, 26, -92, -44, -93, -2, 28, -52, -110, -6, 9, 3, 98, 39, -28, 100, 61, 53, -66, 51, -78, -47, 52, -7, 22, -44, -46, -49, -72, 8, 22, 36, 78, 51, 21, -19, -7, -49, -17, 100, -47, -43, -19, -25, 69, -18, -19, 26, -48, -47, -9, -74, 4, 71, 50, -15, -6, -43, -96, -61, -15, 1, 17, -10, 60, -18, -37, -3, 1, -81, -8, -102, 62, -7),
  48 => (22, -77, 1, -7, 80, 12, 11, -32, 19, 54, 21, 52, 24, -8, 13, -75, -22, 13, 54, -16, -33, -4, 14, 58, 10, 12, 20, -9, 121, 2, -12, 15, 129, 10, 83, 44, -12, 39, 10, 5, -1, 8, 8, 61, -4, -27, 44, -2, -85, 22, -105, 29, 59, 11, -8, 38, -70, -5, -49, 54, -39, -89, -85, -56, 59, -40, 82, -30, -77, 8, 60, 27, -73, 19, 20, -13, -12, 81, 35, 4, 14, -58, -70, 68, -25, 52, 12, -5, 5, -13, 13, 25, 4, -28, -48, -8, -28, 6, 20, 32, 27, 135, 8, -26, -1, -59, 75, 81, 58, 9, 47, -66, -17, -80, 74, 48, -110, 6, 12, -73, 40, 39, -5, -65, 57, 11, 47, -28),
  49 => (70, -44, -58, -19, -73, -43, 29, 5, -2, -23, 36, 15, -51, 45, 63, 50, -58, -94, -10, -3, 2, 0, -9, -35, -31, -28, 4, -25, 44, 4, 61, 84, -110, -46, 8, -20, 42, -57, 11, -3, 37, 29, -32, 105, 58, 22, 96, 47, -17, -7, 114, -12, -28, 30, -67, -33, 34, 7, -59, -41, 31, -42, -63, 16, 10, 7, 44, 84, 55, -40, -69, 46, -19, -73, 75, 30, 23, -41, 115, 66, 17, 4, -57, 23, 52, 38, -10, -12, 27, 20, -50, 20, 23, -9, -72, 31, -34, -79, 69, 91, -75, -90, -20, 16, -17, -32, -22, 23, -62, -67, 23, 26, 85, 75, 2, 49, 55, 86, -60, -38, 57, -28, 51, 33, 13, 27, -29, 2),
  50 => (68, 11, -35, 68, -81, 16, 45, 8, 27, 32, -106, -55, -26, 6, 41, -21, -116, -2, 91, 63, -63, -34, -26, 32, 19, -93, -19, 4, -57, 18, 99, 89, -6, -13, -36, 48, 75, -24, -27, -95, -8, 5, -18, 37, 53, 19, 27, 48, 30, 16, -7, 0, -102, 66, -66, 60, 1, -20, 6, -33, 103, -51, 37, 24, 34, 41, -11, 69, 26, 6, -60, 10, -26, 46, -7, -45, -1, -44, 10, 42, 38, 24, -19, -35, 33, 8, -32, -15, 32, -47, 10, -80, -92, 32, -9, -32, -23, 11, -22, 46, -50, 5, -96, 28, 55, 1, 76, 78, -10, -31, 63, 44, -18, -49, 95, 25, -4, -30, 90, -30, 25, 36, -58, -4, 83, -4, 84, -4),
  51 => (-81, -47, -135, -42, 40, -25, 27, -3, -45, 3, 36, 58, -96, -22, 36, 40, 18, 18, -1, -19, 30, -112, -108, 9, -102, 103, -15, -125, -6, -17, 25, -30, 62, -1, 77, -59, 24, 94, 27, 31, -69, -83, 21, -43, -38, -1, 7, -34, 18, 96, -60, 60, 48, 49, 55, 50, 6, 5, -20, 66, 18, 45, -30, 31, 16, -55, -12, 17, 44, 30, 35, 2, 25, -12, 27, 52, 30, 67, 17, -40, 56, -8, 43, 45, -10, -31, 72, -12, -19, -66, -28, 27, 46, -25, -3, -43, 13, -53, -31, -59, 94, 78, 24, -79, 1, 14, 57, 38, 79, 40, 18, -23, 18, -11, 68, -32, -37, -44, 39, -51, -24, 37, 4, -50, -2, 0, 15, 20),
  52 => (2, 27, 28, -54, -17, 1, 91, 43, -70, 8, 24, 3, 26, -58, 40, -4, 33, 38, 6, -25, -25, 126, 70, 69, 0, 12, -57, 96, 31, -38, -40, 28, 56, 102, 23, 29, -60, -89, 15, 11, -77, 28, -69, -44, 7, -24, -14, 8, -39, -66, 31, -46, 7, -44, -1, -44, -2, 31, 40, 23, 13, -45, -3, -100, 14, 74, -28, -9, -21, -79, -28, 43, -82, -35, -47, 71, -59, 58, -32, -51, 40, -25, 20, 21, 0, -19, -17, -98, -34, 17, 37, -84, 45, 32, -67, -20, 76, 45, 77, -22, -106, 59, 52, 9, 8, 61, 58, 31, 31, 59, 10, 59, -60, -43, -35, -18, 2, -23, 53, 10, -22, 2, -60, -110, 0, -1, -1, 3),
  53 => (27, 94, 91, -39, -77, -54, -54, 16, 19, 12, -47, -105, -31, 24, -64, 12, 40, -45, -72, 24, -29, 121, 40, -5, 43, -12, 101, 87, -23, 43, 21, 1, -82, 29, -43, -71, -69, -16, 39, -58, 52, 29, 53, -15, -11, -87, -24, -28, 109, -19, -12, -40, -92, -11, 7, 4, -22, 59, -34, 12, -35, 62, 42, -33, 18, 69, -42, -30, 7, -11, 28, -50, 1, -39, 1, -68, 20, -95, -17, -29, -30, 51, 38, -52, 34, -1, -88, 8, -63, 12, 54, 0, -12, -26, 79, -17, -7, 33, 5, -61, -77, -58, -5, 88, 22, -40, -18, -57, -8, 66, -12, 5, 19, -25, -15, -12, -52, -49, -33, 91, 31, 30, 0, 4, -3, -109, 1, 20),
  54 => (42, 48, -58, -49, 32, -36, -22, -30, 53, -19, 41, -18, -8, 113, 0, 36, 74, 28, 9, 19, 34, -51, -13, -3, -15, 21, 82, -13, 8, -13, -92, -39, -16, 22, 3, 23, -59, 44, -52, 55, -43, 7, 69, 22, -43, -47, 2, -45, -1, 35, 6, 22, -2, -75, -22, 25, 111, 17, 53, 10, -9, 12, 34, 93, -5, -5, -17, -47, 70, 53, 29, 74, 34, 16, 76, 2, -65, -25, -60, -29, -26, 13, 11, 28, -25, -72, 13, -69, 30, -22, 0, 69, -71, -3, 9, 54, 19, -5, 26, 26, 43, -58, -29, 70, 22, -29, -57, 2, -14, 58, -31, 50, 42, 67, 15, 20, 109, 80, 52, 38, 64, -10, -15, 87, -53, 151, -43, -37),
  55 => (-53, 1, -85, -23, -14, -2, 30, -41, 63, 34, -8, 44, -98, -89, -41, 93, -2, 57, -45, 87, 11, -48, 3, 7, -53, 16, 64, -21, -102, -37, 15, -61, 6, 1, 10, -63, -82, 24, 84, 12, 12, -3, 26, -37, 13, 55, -77, -33, 16, 88, 25, 86, -48, 37, 40, 67, 61, 5, -27, 13, -10, -3, 27, 27, -52, -44, -10, 27, 42, 2, 36, -32, 3, 71, 0, 42, -3, 4, 2, -75, -9, 11, 35, 9, 58, 31, 48, 17, 16, 33, -9, -4, -17, 49, 72, -138, 90, -46, -28, 36, 43, 23, 7, 41, 61, 6, 11, 77, -16, 52, -30, 44, 23, 28, 41, -91, -52, 13, 77, -33, -12, 59, -10, 25, 48, -34, -30, 68),
  56 => (-145, 10, -77, 46, 117, 54, 25, -43, 40, -5, 44, 56, -46, -102, 16, -12, 4, 23, 11, 26, 58, -40, -10, 8, -34, 65, 15, 17, -30, -82, 42, -35, 51, 19, 41, -79, 10, 6, 36, 58, -22, -135, -29, -148, -2, 44, -95, -44, 27, 28, -14, 50, 47, -12, -5, 35, 26, -18, 0, -9, -6, -3, 50, 30, -77, -56, 47, 51, -38, 33, 10, 41, -14, 72, -71, 9, 64, 87, 27, -131, -7, -17, 23, 10, 11, 20, 47, 45, 3, 13, -43, -14, 0, 20, 19, -154, 1, -44, 5, -40, 26, 92, 30, 1, -42, 60, 40, 34, 27, 47, -9, 9, -50, 21, -33, -74, -22, -29, 54, 24, -155, 38, 22, -40, 33, -18, 19, 78),
  57 => (22, -36, 18, 33, 73, -50, -8, -5, 26, -41, 72, 45, 57, 67, 18, 27, 61, 7, -46, -83, 70, 6, -42, -28, 30, -39, 24, -61, 84, -15, -13, 21, 8, 61, 101, -19, 38, 47, -8, 92, -52, 77, 26, 38, 26, -41, -38, 8, 2, 20, 26, 0, 124, -20, 30, -67, -37, 21, -58, -21, -22, 92, -116, -36, -14, -43, 74, 23, -11, 21, 33, 6, -64, -3, 72, 39, -30, 77, -63, -23, -70, -77, 0, 8, -15, -24, 8, -14, -55, -32, -22, 34, 57, -63, -74, 62, -30, 45, 19, -80, 37, 20, 62, 10, -41, 42, -52, -21, -17, -37, -101, 23, 26, -12, -11, 26, -36, 3, -32, -8, 7, -25, -28, 8, -55, 16, -42, -84),
  58 => (-51, 42, -42, 60, 69, -32, 70, 29, 6, -67, 34, -63, -39, 48, 79, 4, 79, 17, -8, -1, 31, 30, 20, -62, 20, -20, 33, 22, 62, -117, 0, 51, -40, 130, -22, 22, 35, -35, -74, 56, -37, 0, 29, -113, -13, -21, -61, -53, -57, -13, 19, -7, 55, -28, -7, -93, -16, 51, 6, -16, 41, 66, -24, -51, -50, 39, 15, 25, 16, 33, 6, 76, -81, -38, -10, -55, -46, -23, -38, -46, -35, -41, 29, -14, -17, -18, 39, -25, -1, 23, 25, 2, -7, 20, -41, -26, 84, 28, 73, -39, -57, -26, 57, 14, 23, -31, -5, -24, 16, 78, -39, 37, -87, 47, -40, -41, 34, 32, 49, -16, -77, 34, -45, -10, -85, -17, 24, -63),
  59 => (44, 21, 63, 52, -6, 1, -57, -91, 27, 14, -59, 17, 140, -27, 9, 39, 24, 55, 32, -53, -25, 77, 44, 35, 37, -63, 17, 16, 16, -18, 6, -7, 17, 70, 25, 28, 56, 11, 32, -54, -10, -23, -49, 25, -38, 22, -3, 102, -4, -42, 21, -91, 18, 44, 52, -37, -110, 36, -69, -27, -44, 90, 80, -79, -64, 75, 13, 34, 33, -23, 15, -10, 78, 73, -41, -26, -77, 0, -11, 50, 23, -91, -20, 0, -28, -29, -52, 28, 69, -60, 70, 2, -21, -43, -24, -25, 63, 44, -48, -25, -69, 34, 19, 12, -68, 63, 55, 5, 43, 89, -19, -16, -38, 3, 39, -3, 5, 36, 21, -4, 7, 91, -10, 94, 16, -27, -59, -96),
  60 => (-64, 22, 36, 47, 29, 38, 77, 2, 85, -50, 40, 74, 31, 4, 83, -37, 6, 34, 25, -74, -1, 52, -12, 19, 49, 12, 50, -10, -23, -29, 2, -90, -36, -37, -16, 0, -4, 87, -91, 1, -152, -52, 70, -42, -80, 51, -77, -75, 44, -15, 43, -87, 11, 1, -54, -27, 67, -51, 70, -42, 80, 63, 92, -51, -43, -15, 64, -26, 9, -20, 12, 34, -2, -24, 26, -10, -19, 13, -43, -85, -45, 24, 25, -95, -30, -59, -33, 21, -60, -49, 29, -28, -22, 48, 6, -13, 44, 27, -36, 3, 26, -14, -71, 52, -21, 29, -16, 42, -25, 3, 31, -12, 61, 19, 26, 23, 19, 55, -38, 67, -13, 8, 87, 36, -63, 57, 108, 85),
  61 => (57, -5, 38, -45, -40, -37, -116, 19, -82, 1, -1, -27, 18, 13, -80, 19, -29, -122, 38, -9, -29, 94, 10, -18, 47, -26, -44, 18, 21, 3, -60, -52, 43, -29, 21, -24, -13, -86, -34, 51, -7, 74, 38, 46, 7, -46, 31, 27, 58, 5, -48, 1, -5, -69, -16, 62, -6, -16, 2, 2, -20, -12, -5, -11, 56, -19, -38, -33, -127, -43, 29, -37, -18, 10, 50, 15, -39, 21, -11, 42, 16, -35, 51, -32, 14, 7, 58, -75, -15, -53, 25, -27, 37, -56, 27, 78, -35, 6, -46, -40, -24, 47, -5, 26, -31, -31, 24, 35, 22, 37, 102, 32, -7, -122, 64, 43, -133, -59, 17, 2, 101, 30, -144, -59, 95, 15, -56, -8),
  62 => (-84, -14, -11, -15, 41, -34, 4, -24, -54, -3, 48, 76, -10, -44, -16, 1, -12, -59, -1, -51, 17, -5, 0, 23, -2, 65, -53, 16, 61, -96, -34, -44, 116, 4, 86, -23, 19, -58, 78, 24, 43, 39, -98, -46, -15, -11, 56, 26, -1, 49, -15, 68, 30, -94, 13, 54, -44, 23, -54, -17, 30, 23, 32, -17, 49, -34, 8, -4, -16, 59, -16, -65, -10, 66, -29, 68, 18, 105, -40, 12, 78, -78, -13, -21, -25, 44, -68, -47, -4, 21, -41, -43, 42, 4, 33, -83, 0, -40, 47, 61, -8, 135, 54, -26, -26, 39, 98, -23, 83, -41, 7, 15, -33, -41, -60, -33, -113, -34, -45, -71, -87, 23, -51, 19, 146, -65, -80, -1),
  63 => (-5, -72, 73, 65, -8, 35, -27, 68, 163, -13, 0, -39, 76, -8, -40, -14, -6, 91, 26, 67, 39, 51, 65, -11, 60, -28, 17, 68, -72, 22, -23, 1, 10, 65, 43, -24, -44, 62, -35, -5, -14, -57, 13, -9, -18, 52, -40, 31, 30, -97, -8, -57, 28, -21, 5, 43, -1, 40, -7, -33, 23, -52, 92, -79, -24, -5, 10, -53, 3, -48, -19, -66, 24, 26, -59, -4, -12, 55, -43, -31, -22, 18, 40, -31, -86, -18, -64, 46, 51, -23, 129, -9, -31, -9, 8, -67, -13, 88, -69, 38, 10, 40, -57, 9, 87, 86, 30, 42, 31, -8, 73, 11, 0, -69, 27, -51, -72, -17, -19, -47, 10, 67, 52, 48, 72, 23, 67, 69)
);


constant weight_matrix_layer6 :  weight_matrix_layer6_type := (
  0 => (40, 2, -129, 44, -106, 61, -43, 70, -76, -111, -62, 54, -70, -92, -68, 52, -84, -124, 23, 19, 23, 72, 12, -49, 51, 67, -41, -64, -109, 57, -37, 28, 11, 63, 0, -66, -110, 81, -95, 9, 68, 61, -70, 43, 75, -126, -41, 33, 3, -35, -134, 81, 57, -124, -88, 67, 89, 38, 63, 11, -120, -81, 61, -138),
  1 => (-126, 64, 47, -57, 92, -40, -140, 32, -56, -28, -30, 81, -121, 104, 84, -59, -138, 4, -156, -136, 98, -53, -78, -65, -22, -121, 82, -187, 73, 10, -129, -60, -103, -63, 30, 57, 77, 46, -57, -115, 38, 44, -28, 32, 81, -48, -55, -24, 70, -121, -33, 75, -75, -115, 82, -42, -71, 79, -76, -129, -88, 53, 54, -104),
  2 => (-79, 13, 81, -64, -65, 87, 51, -87, -126, -126, 55, 46, 55, -25, 102, 52, -35, -100, 52, 50, 62, 28, -75, 64, 70, 74, -43, -78, 77, -139, 46, -12, 63, -42, 11, -91, 62, -42, 52, -10, -130, -108, -63, 86, -77, -81, -104, -63, -95, 2, -85, -12, 79, 68, 79, 34, -137, 5, 47, 59, 0, -46, -35, 78),
  3 => (86, 109, -75, -121, 54, 59, -145, -100, 37, 61, -128, 60, 78, 21, -68, 40, 82, -43, 27, 68, -102, -125, -81, 48, -72, -89, 40, 42, -100, -114, 55, 80, 70, 40, 52, -58, 69, 43, 53, -131, -54, -143, -15, 31, 54, -20, 20, -122, -37, -2, 55, -109, -4, 82, -50, 22, -113, -78, -82, 45, -145, 52, 56, -106),
  4 => (-148, -86, 86, 44, -111, -40, 67, -129, -108, -37, 53, -86, -81, 81, 78, -133, -84, -82, -15, -62, 75, 57, -12, 71, -76, 81, 35, 49, 73, 46, -77, -98, -50, 18, -35, 62, -113, -111, -130, 63, -35, 63, 55, 66, 34, -75, -144, -110, -38, 76, 28, 45, -61, -133, 62, 66, 52, -95, -95, -104, 76, -38, 55, 88),
  5 => (71, 65, 17, 55, 39, -24, -121, 44, -47, 72, -97, 69, 78, -89, -16, 37, 80, 78, -1, 67, -110, -123, 78, -51, 47, 53, -156, 36, 14, 43, 19, 81, -77, 76, -132, -95, -74, -47, 5, -119, 55, 60, -50, -3, -72, 72, -88, 18, -98, -144, 27, -121, 19, 73, 64, -26, 45, 10, 71, 63, 52, 25, -107, 5),
  6 => (-12, 37, -115, 65, 14, -118, 44, 94, -52, 21, 53, 10, -66, -24, -76, 23, 53, 43, -35, -63, 97, 41, -15, 64, 67, 62, 43, -82, 68, 43, -22, 71, -31, -120, 80, -142, -101, 49, -111, 67, 57, 75, -132, -66, -60, -54, 47, -83, -121, 63, -140, -20, -66, -6, 72, -84, -39, 58, 12, -82, 87, -103, -151, 26),
  7 => (-107, -92, 38, -108, 56, 52, 40, 45, 30, -83, -1, -165, 83, 81, -10, -190, -38, 46, -146, 72, 12, -26, -137, -72, 101, -75, 34, -97, 14, -146, -116, -98, 10, -56, 55, 48, 59, 52, 56, -62, 57, -116, 74, -77, -41, 37, 41, -6, 48, -49, 81, -60, 79, 17, -119, -102, -58, 41, -173, 91, -76, 57, 55, 23),
  8 => (-2, -43, -149, 79, -36, -56, 38, 58, 40, 96, -113, -10, -98, -138, 28, -57, -74, -113, 23, 39, -39, -28, -89, -73, -57, 63, -86, 70, -137, -71, 58, -51, 70, 80, 13, -105, -55, 66, 61, 43, 60, -74, 36, -99, -68, -55, 52, 62, -50, 54, 65, -97, -117, -72, -37, -44, 8, -23, 28, -60, -106, -152, -99, -108),
  9 => (39, -29, 55, -59, 13, -8, 28, -60, 54, 74, -99, -109, 40, -30, 25, -124, -95, -66, -183, -73, -109, -21, -5, 14, -80, -138, -123, 49, -132, 35, -22, -39, -144, 82, -85, 43, -63, 57, 67, -25, -118, 59, 61, -18, 98, 84, 50, 54, 50, -104, 47, 51, -89, 0, -84, 47, 76, -138, -81, 4, 64, -81, 54, 48)
);

end package Layer4_6_Weights;

package body Layer4_6_Weights is
end package body;